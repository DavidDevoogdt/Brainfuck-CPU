* NGSPICE file created from BFCPU.ext - technology: scmos

.global Vdd Gnd 

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

.subckt BFCPU vdd gnd clk INPD<0> INPD<1> INPD<2> INPD<3> INPD<4> INPD<5> INPD<6>
+ INPD<7> INPD<8> INPD<9> INPD<10> INPD<11> INPD<12> INPD<13> INPD<14> INPD<15> RDATA<0>
+ RDATA<1> RDATA<2> RDATA<3> RDATA<4> RDATA<5> RDATA<6> RDATA<7> RF WF NEXTOP<0> NEXTOP<1>
+ NEXTOP<2> IR OW OUTPD<0> OUTPD<1> OUTPD<2> OUTPD<3> OUTPD<4> OUTPD<5> OUTPD<6> OUTPD<7>
+ OUTPD<8> OUTPD<9> OUTPD<10> OUTPD<11> OUTPD<12> OUTPD<13> OUTPD<14> OUTPD<15> reset
+ RD WD WDATA<0> WDATA<1> WDATA<2> WDATA<3> WDATA<4> WDATA<5> WDATA<6> WDATA<7> DP<0>
+ DP<1> DP<2> DP<3> DP<4> DP<5> DP<6> DP<7> DP<8> DP<9> DP<10> DP<11> DP<12> DP<13>
+ DP<14> PCDELTA<0> PCDELTA<1> PCDELTA<2> PCDELTA<3> PCDELTA<4> PCDELTA<5> PCDELTA<6>
+ PCDELTA<7> PCDELTA<8> PCDELTA<9> PCDELTA<10> PCDELTA<11> PCDELTA<12> PCDELTA<13>
+ PCDELTA<14> PCDELTA<15>
XFILL_1_2 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XNAND2X1_16 INVX2_3/A RDATA<5> gnd NAND2X1_16/Y vdd NAND2X1
XBUFX2_42 BUFX2_68/A gnd PCDELTA<8> vdd BUFX2
XBUFX2_43 BUFX2_68/A gnd PCDELTA<9> vdd BUFX2
XBUFX2_40 BUFX2_68/A gnd PCDELTA<6> vdd BUFX2
XBUFX2_68 BUFX2_68/A gnd BUFX2_68/Y vdd BUFX2
XBUFX2_33 XOR2X1_1/B gnd OW vdd BUFX2
XXOR2X1_1 XOR2X1_1/A XOR2X1_1/B gnd XOR2X1_1/Y vdd XOR2X1
XBUFX2_30 BUFX2_30/A gnd OUTPD<13> vdd BUFX2
XBUFX2_67 BUFX2_38/A gnd BUFX2_67/Y vdd BUFX2
XBUFX2_46 BUFX2_38/A gnd PCDELTA<12> vdd BUFX2
XBUFX2_72 BUFX2_38/A gnd BUFX2_72/Y vdd BUFX2
XBUFX2_66 BUFX2_38/A gnd BUFX2_66/Y vdd BUFX2
XBUFX2_38 BUFX2_38/A gnd PCDELTA<4> vdd BUFX2
XBUFX2_32 BUFX2_32/A gnd OUTPD<15> vdd BUFX2
XDFFPOSX1_9 BUFX2_24/A BUFX4_10/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XFILL_0_1_1 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XBUFX2_24 BUFX2_24/A gnd OUTPD<7> vdd BUFX2
XBUFX2_17 BUFX2_17/A gnd OUTPD<0> vdd BUFX2
XDFFPOSX1_2 BUFX2_17/A BUFX4_10/Y AOI21X1_7/Y gnd vdd DFFPOSX1
XBUFX2_51 BUFX2_51/A gnd WD vdd BUFX2
XBUFX2_50 BUFX2_50/A gnd RD vdd BUFX2
XDFFPOSX1_45 INVX1_2/A BUFX4_10/Y NAND3X1_23/Y gnd vdd DFFPOSX1
XNAND3X1_23 NAND2X1_41/Y OAI21X1_55/Y NOR3X1_19/Y gnd NAND3X1_23/Y vdd NAND3X1
XBUFX2_34 BUFX2_34/A gnd PCDELTA<0> vdd BUFX2
XNAND2X1_41 INVX1_35/Y OAI21X1_53/Y gnd NAND2X1_41/Y vdd NAND2X1
XOAI21X1_55 NOR3X1_13/Y OAI21X1_54/Y NEXTOP<2> gnd OAI21X1_55/Y vdd OAI21X1
XNOR3X1_16 INVX1_37/A NOR2X1_53/Y NOR3X1_16/C gnd NOR3X1_16/Y vdd NOR3X1
XOAI21X1_54 INVX4_3/Y NOR3X1_9/B OAI22X1_3/C gnd OAI21X1_54/Y vdd OAI21X1
XFILL_0_0_1 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XNOR2X1_53 NOR3X1_9/B NOR2X1_53/B gnd NOR2X1_53/Y vdd NOR2X1
XNAND3X1_15 RF INVX2_11/Y INVX4_3/Y gnd NOR2X1_53/B vdd NAND3X1
XNOR3X1_11 NEXTOP<0> NOR3X1_11/B INVX1_30/A gnd NOR3X1_11/Y vdd NOR3X1
XOAI21X1_52 OAI21X1_52/A NOR3X1_11/B INVX2_11/Y gnd OAI21X1_53/C vdd OAI21X1
XOAI21X1_53 NOR3X1_11/Y INVX2_11/Y OAI21X1_53/C gnd OAI21X1_53/Y vdd OAI21X1
XINVX2_11 BUFX4_1/Y gnd INVX2_11/Y vdd INVX2
XNOR3X1_13 NOR3X1_9/A INVX2_12/Y NOR3X1_9/B gnd NOR3X1_13/Y vdd NOR3X1
XNOR2X1_46 NEXTOP<0> INVX2_12/Y gnd NOR3X1_9/C vdd NOR2X1
XNOR3X1_9 NOR3X1_9/A NOR3X1_9/B NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XNAND2X1_35 BUFX4_1/Y INVX4_3/Y gnd NOR3X1_9/A vdd NAND2X1
XNOR2X1_56 NOR3X1_9/A NOR3X1_9/B gnd NOR2X1_56/Y vdd NOR2X1
XAOI21X1_24 INVX2_12/Y NOR2X1_56/Y AOI21X1_24/C gnd AOI21X1_24/Y vdd AOI21X1
XINVX2_12 WF gnd INVX2_12/Y vdd INVX2
XBUFX2_60 BUFX2_60/A gnd reset vdd BUFX2
XFILL_2_1 gnd vdd FILL
XBUFX4_21 BUFX4_22/A gnd BUFX2_68/A vdd BUFX4
XDFFPOSX1_27 XOR2X1_1/B BUFX4_10/Y XOR2X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_15 BUFX2_30/A BUFX4_10/Y NOR2X1_30/Y gnd vdd DFFPOSX1
XINVX1_18 BUFX2_30/A gnd INVX1_18/Y vdd INVX1
XNOR2X1_30 INVX1_18/Y BUFX4_16/Y gnd NOR2X1_30/Y vdd NOR2X1
XBUFX4_22 BUFX4_22/A gnd BUFX2_38/A vdd BUFX4
XBUFX4_13 BUFX4_16/A gnd XOR2X1_1/A vdd BUFX4
XBUFX4_16 BUFX4_16/A gnd BUFX4_16/Y vdd BUFX4
XAOI21X1_14 INVX2_2/Y BUFX4_16/Y NOR2X1_24/Y gnd DFFPOSX1_9/D vdd AOI21X1
XNOR2X1_24 BUFX2_24/A BUFX4_16/Y gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_17 BUFX2_17/A BUFX4_16/Y gnd AOI21X1_7/C vdd NOR2X1
XAOI21X1_7 INVX2_5/Y BUFX4_16/Y AOI21X1_7/C gnd AOI21X1_7/Y vdd AOI21X1
XFILL_1_1_1 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XNAND2X1_4 INVX1_1/A INVX1_2/A gnd NOR2X1_5/A vdd NAND2X1
XNOR2X1_6 NOR2X1_5/A NOR2X1_6/B gnd BUFX2_51/A vdd NOR2X1
XNOR2X1_5 NOR2X1_5/A OR2X2_1/Y gnd BUFX2_50/A vdd NOR2X1
XNOR3X1_17 NOR3X1_15/C NOR3X1_15/B NOR2X1_54/Y gnd NOR3X1_19/A vdd NOR3X1
XNOR3X1_15 NOR3X1_15/A NOR3X1_15/B NOR3X1_15/C gnd NOR3X1_16/C vdd NOR3X1
XNOR3X1_19 NOR3X1_19/A NOR3X1_19/B OAI22X1_3/Y gnd NOR3X1_19/Y vdd NOR3X1
XNAND2X1_40 NEXTOP<1> INVX1_33/Y gnd NOR3X1_15/A vdd NAND2X1
XINVX1_33 NEXTOP<2> gnd INVX1_33/Y vdd INVX1
XNOR2X1_54 NEXTOP<2> INVX2_13/Y gnd NOR2X1_54/Y vdd NOR2X1
XNAND2X1_44 INVX1_31/A NOR2X1_42/Y gnd NAND3X1_25/A vdd NAND2X1
XNOR2X1_52 INVX1_35/Y NOR2X1_52/B gnd NOR2X1_52/Y vdd NOR2X1
XAOI21X1_23 INVX2_13/Y INVX4_4/Y OAI22X1_3/C gnd NOR2X1_52/B vdd AOI21X1
XINVX2_13 NEXTOP<1> gnd INVX2_13/Y vdd INVX2
XOAI21X1_48 INVX1_33/Y NEXTOP<0> INVX2_13/Y gnd NOR2X1_48/A vdd OAI21X1
XOAI22X1_3 OAI22X1_3/A NOR2X1_44/A OAI22X1_3/C INVX4_4/Y gnd OAI22X1_3/Y vdd OAI22X1
XFILL_1_0_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XNOR2X1_43 NEXTOP<2> NEXTOP<1> gnd NOR2X1_44/A vdd NOR2X1
XNAND3X1_22 NEXTOP<2> NEXTOP<1> NEXTOP<0> gnd OAI21X1_52/A vdd NAND3X1
XNAND2X1_31 NEXTOP<2> NEXTOP<1> gnd INVX1_30/A vdd NAND2X1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XNOR2X1_44 NOR2X1_44/A INVX1_30/Y gnd INVX1_31/A vdd NOR2X1
XOAI21X1_56 INVX1_30/Y NOR2X1_44/A NOR2X1_42/Y gnd NAND3X1_24/A vdd OAI21X1
XNAND2X1_42 INVX4_3/Y NOR2X1_47/Y gnd OAI22X1_3/A vdd NAND2X1
XNOR2X1_47 INVX1_1/A INVX1_2/A gnd NOR2X1_47/Y vdd NOR2X1
XNAND3X1_16 NEXTOP<0> INVX4_3/Y NOR2X1_47/Y gnd NOR2X1_48/B vdd NAND3X1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XNAND3X1_24 NAND3X1_24/A AOI21X1_24/Y NOR3X1_20/Y gnd NAND3X1_24/Y vdd NAND3X1
XDFFPOSX1_46 INVX1_1/A BUFX4_8/Y NAND3X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_1 BUFX2_60/A BUFX4_8/Y vdd gnd vdd DFFPOSX1
XFILL_3_1 gnd vdd FILL
XBUFX2_23 BUFX2_23/A gnd OUTPD<6> vdd BUFX2
XDFFPOSX1_5 BUFX2_20/A BUFX4_10/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XNOR2X1_22 BUFX2_22/A XOR2X1_1/A gnd NOR2X1_22/Y vdd NOR2X1
XAOI21X1_12 INVX2_1/Y XOR2X1_1/A NOR2X1_22/Y gnd DFFPOSX1_7/D vdd AOI21X1
XNOR2X1_23 BUFX2_23/A XOR2X1_1/A gnd NOR2X1_23/Y vdd NOR2X1
XDFFPOSX1_8 BUFX2_23/A BUFX4_7/Y DFFPOSX1_8/D gnd vdd DFFPOSX1
XNOR2X1_32 INVX1_20/Y XOR2X1_1/A gnd NOR2X1_32/Y vdd NOR2X1
XINVX1_20 BUFX2_32/A gnd INVX1_20/Y vdd INVX1
XDFFPOSX1_17 BUFX2_32/A BUFX4_7/Y NOR2X1_32/Y gnd vdd DFFPOSX1
XBUFX2_52 INVX2_5/A gnd WDATA<0> vdd BUFX2
XBUFX2_26 BUFX2_26/A gnd OUTPD<9> vdd BUFX2
XFILL_2_1_1 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XDFFPOSX1_11 BUFX2_26/A BUFX4_7/Y NOR2X1_26/Y gnd vdd DFFPOSX1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XNAND2X1_39 INVX1_1/A NOR3X1_15/B gnd INVX1_35/A vdd NAND2X1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XAND2X2_15 INVX1_2/A INVX4_3/A gnd NOR3X1_15/B vdd AND2X2
XNOR2X1_42 NOR3X1_15/B NOR3X1_15/C gnd NOR2X1_42/Y vdd NOR2X1
XOAI21X1_46 INVX1_2/A INVX4_3/A INVX2_10/Y gnd NOR3X1_15/C vdd OAI21X1
XINVX2_10 INVX1_1/A gnd INVX2_10/Y vdd INVX2
XNOR3X1_18 OR2X2_4/A NOR3X1_18/B NOR2X1_55/Y gnd NOR3X1_19/B vdd NOR3X1
XNAND3X1_25 NAND3X1_25/A NOR2X1_60/Y NAND3X1_25/C gnd BUFX2_34/A vdd NAND3X1
XNOR2X1_55 NEXTOP<2> INVX4_4/Y gnd NOR2X1_55/Y vdd NOR2X1
XOAI21X1_51 NOR3X1_13/Y OAI21X1_51/B NEXTOP<1> gnd NAND3X1_21/B vdd OAI21X1
XNAND3X1_21 NOR2X1_52/Y NAND3X1_21/B NOR3X1_16/Y gnd NAND3X1_21/Y vdd NAND3X1
XNOR2X1_60 NOR3X1_13/Y OAI22X1_4/Y gnd NOR2X1_60/Y vdd NOR2X1
XOAI22X1_4 INVX2_10/Y INVX4_3/Y OAI22X1_3/A NOR2X1_48/A gnd OAI22X1_4/Y vdd OAI22X1
XFILL_2_0_1 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XNOR2X1_57 INVX4_4/Y OAI22X1_3/C gnd NOR3X1_20/C vdd NOR2X1
XOAI22X1_2 NOR3X1_9/B NOR2X1_53/B OAI22X1_3/C OAI22X1_2/D gnd NOR3X1_10/C vdd OAI22X1
XAOI21X1_25 NEXTOP<2> INVX1_34/Y NEXTOP<1> gnd NOR2X1_58/A vdd AOI21X1
XNOR2X1_58 NOR2X1_58/A OAI22X1_3/A gnd NOR3X1_20/A vdd NOR2X1
XNOR3X1_20 NOR3X1_20/A INVX1_37/A NOR3X1_20/C gnd NOR3X1_20/Y vdd NOR3X1
XNOR2X1_48 NOR2X1_48/A NOR2X1_48/B gnd NOR3X1_10/A vdd NOR2X1
XOAI21X1_47 INVX1_31/Y NEXTOP<0> NOR2X1_42/Y gnd OAI21X1_47/Y vdd OAI21X1
XNOR3X1_10 NOR3X1_10/A NOR3X1_9/Y NOR3X1_10/C gnd NOR3X1_10/Y vdd NOR3X1
XNAND2X1_43 INVX1_1/A INVX4_3/Y gnd OAI21X1_57/A vdd NAND2X1
XOAI21X1_57 OAI21X1_57/A BUFX4_1/Y OR2X2_4/B gnd AOI21X1_24/C vdd OAI21X1
XDFFPOSX1_44 INVX4_3/A BUFX4_8/Y NAND3X1_21/Y gnd vdd DFFPOSX1
XFILL_4_3 gnd vdd FILL
XFILL_4_2 gnd vdd FILL
XFILL_4_1 gnd vdd FILL
XBUFX2_41 BUFX2_68/A gnd PCDELTA<7> vdd BUFX2
XBUFX2_20 BUFX2_20/A gnd OUTPD<3> vdd BUFX2
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XNOR2X1_20 BUFX2_20/A BUFX4_15/Y gnd NOR2X1_20/Y vdd NOR2X1
XAOI21X1_10 INVX1_6/Y BUFX4_15/Y NOR2X1_20/Y gnd DFFPOSX1_5/D vdd AOI21X1
XDFFPOSX1_7 BUFX2_22/A BUFX4_10/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XAOI21X1_13 INVX4_2/Y BUFX4_15/Y NOR2X1_23/Y gnd DFFPOSX1_8/D vdd AOI21X1
XDFFPOSX1_21 INVX1_6/A BUFX4_10/Y OAI21X1_10/Y gnd vdd DFFPOSX1
XOAI21X1_10 AND2X2_4/Y OAI21X1_7/Y OAI21X1_9/Y gnd OAI21X1_10/Y vdd OAI21X1
XAND2X2_4 AND2X2_4/A INVX1_6/A gnd AND2X2_4/Y vdd AND2X2
XOAI21X1_7 AND2X2_4/A INVX1_6/A NOR2X1_2/Y gnd OAI21X1_7/Y vdd OAI21X1
XBUFX4_10 clk gnd BUFX4_10/Y vdd BUFX4
XFILL_3_1_1 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XBUFX4_7 clk gnd BUFX4_7/Y vdd BUFX4
XINVX1_14 BUFX2_26/A gnd INVX1_14/Y vdd INVX1
XNOR2X1_26 INVX1_14/Y BUFX4_17/Y gnd NOR2X1_26/Y vdd NOR2X1
XNOR2X1_45 INVX1_1/A BUFX4_1/Y gnd NOR2X1_45/Y vdd NOR2X1
XNAND2X1_33 NOR2X1_45/Y NOR3X1_15/B gnd OAI22X1_3/C vdd NAND2X1
XNOR2X1_59 INVX4_4/A OAI22X1_3/C gnd NOR2X1_59/Y vdd NOR2X1
XAOI21X1_26 INVX4_4/A INVX1_36/Y NOR2X1_59/Y gnd NAND3X1_25/C vdd AOI21X1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XNAND3X1_18 INVX2_10/Y BUFX4_1/Y NOR3X1_15/B gnd INVX1_36/A vdd NAND3X1
XNAND2X1_38 INVX1_2/A INVX2_10/Y gnd NOR3X1_18/B vdd NAND2X1
XNOR3X1_14 INVX4_4/A OR2X2_4/A NOR3X1_18/B gnd INVX1_37/A vdd NOR3X1
XNAND2X1_36 BUFX4_1/Y INVX4_3/A gnd OR2X2_4/A vdd NAND2X1
XINVX4_4 INVX4_4/A gnd INVX4_4/Y vdd INVX4
XOAI21X1_50 NOR3X1_18/B OR2X2_4/A NOR2X1_51/B gnd OAI21X1_51/B vdd OAI21X1
XNOR2X1_50 NEXTOP<0> INVX4_4/Y gnd NOR2X1_50/Y vdd NOR2X1
XOAI21X1_49 INVX1_36/A NOR2X1_50/Y OAI21X1_49/C gnd NOR3X1_12/C vdd OAI21X1
XOAI21X1_59 INVX4_4/Y OAI22X1_3/C INVX1_37/Y gnd OAI21X1_59/Y vdd OAI21X1
XFILL_3_0_1 gnd vdd FILL
XFILL_3_0_0 gnd vdd FILL
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XNAND2X1_34 NEXTOP<0> INVX4_4/Y gnd OAI22X1_2/D vdd NAND2X1
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XOAI21X1_58 NOR3X1_11/Y OR2X2_4/Y INVX1_37/Y gnd BUFX4_22/A vdd OAI21X1
XINVX1_34 NEXTOP<0> gnd INVX1_34/Y vdd INVX1
XNOR2X1_51 INVX1_34/Y NOR2X1_51/B gnd NOR3X1_12/B vdd NOR2X1
XNOR2X1_49 NOR3X1_11/Y OR2X2_4/Y gnd NOR3X1_12/A vdd NOR2X1
XNOR3X1_12 NOR3X1_12/A NOR3X1_12/B NOR3X1_12/C gnd NOR3X1_12/Y vdd NOR3X1
XNAND3X1_20 OAI21X1_47/Y NOR3X1_10/Y NOR3X1_12/Y gnd NAND3X1_20/Y vdd NAND3X1
XNAND2X1_32 INVX1_1/A INVX1_32/Y gnd NOR3X1_9/B vdd NAND2X1
XNAND2X1_37 INVX1_1/A INVX1_2/A gnd OR2X2_4/B vdd NAND2X1
XNOR2X1_25 INVX1_13/Y BUFX4_17/Y gnd NOR2X1_25/Y vdd NOR2X1
XINVX1_13 BUFX2_25/A gnd INVX1_13/Y vdd INVX1
XDFFPOSX1_10 BUFX2_25/A BUFX4_8/Y NOR2X1_25/Y gnd vdd DFFPOSX1
XBUFX2_25 BUFX2_25/A gnd OUTPD<8> vdd BUFX2
XFILL_5_2 gnd vdd FILL
XFILL_5_1 gnd vdd FILL
XINVX1_10 INPD<5> gnd INVX1_10/Y vdd INVX1
XBUFX2_62 BUFX2_68/A gnd BUFX2_62/Y vdd BUFX2
XBUFX2_21 BUFX2_21/A gnd OUTPD<4> vdd BUFX2
XOAI21X1_8 INVX1_6/Y INVX2_3/A OAI21X1_8/C gnd OAI21X1_9/A vdd OAI21X1
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XOAI21X1_9 OAI21X1_9/A INVX2_4/A OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XNOR2X1_21 BUFX2_21/A BUFX4_15/Y gnd NOR2X1_21/Y vdd NOR2X1
XAOI21X1_11 INVX2_6/Y BUFX4_15/Y NOR2X1_21/Y gnd DFFPOSX1_6/D vdd AOI21X1
XDFFPOSX1_6 BUFX2_21/A BUFX4_7/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XBUFX4_15 BUFX4_16/A gnd BUFX4_15/Y vdd BUFX4
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XDFFPOSX1_18 INVX2_5/A BUFX4_7/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XNOR2X1_11 INVX2_4/A NOR2X1_2/Y gnd INVX1_4/A vdd NOR2X1
XFILL_4_1_1 gnd vdd FILL
XFILL_4_1_0 gnd vdd FILL
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XOAI21X1_2 INVX1_4/Y OAI21X1_1/Y AOI22X1_1/Y gnd OAI21X1_2/Y vdd OAI21X1
XAOI22X1_1 INVX2_5/Y NOR2X1_2/Y XOR2X1_2/A INPD<0> gnd AOI22X1_1/Y vdd AOI22X1
XOAI21X1_1 INVX2_3/Y RDATA<0> NAND2X1_7/Y gnd OAI21X1_1/Y vdd OAI21X1
XNAND2X1_7 INVX2_5/Y INVX2_3/Y gnd NAND2X1_7/Y vdd NAND2X1
XNOR2X1_12 NOR2X1_12/A INVX1_4/Y gnd BUFX4_16/A vdd NOR2X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XNAND2X1_6 NOR2X1_1/Y INVX2_3/Y gnd NOR2X1_12/A vdd NAND2X1
XNOR2X1_1 OR2X2_1/Y NOR2X1_7/A gnd NOR2X1_1/Y vdd NOR2X1
XNOR2X1_7 NOR2X1_7/A NOR2X1_6/B gnd INVX2_4/A vdd NOR2X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XNAND2X1_1 INVX1_2/A INVX1_1/Y gnd NOR2X1_7/A vdd NAND2X1
XOR2X2_1 INVX4_3/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XNAND2X1_5 OR2X2_1/B INVX1_3/Y gnd NOR2X1_6/B vdd NAND2X1
XINVX1_3 INVX4_3/A gnd INVX1_3/Y vdd INVX1
XBUFX2_5 BUFX2_5/A gnd DP<4> vdd BUFX2
XBUFX2_6 BUFX2_6/A gnd DP<5> vdd BUFX2
XDFFPOSX1_32 BUFX2_5/A BUFX4_7/Y XNOR2X1_5/Y gnd vdd DFFPOSX1
XFILL_4_0_1 gnd vdd FILL
XFILL_4_0_0 gnd vdd FILL
XDFFPOSX1_33 BUFX2_6/A BUFX4_7/Y XNOR2X1_6/Y gnd vdd DFFPOSX1
XNAND3X1_17 BUFX4_1/Y INVX4_3/Y AND2X2_16/Y gnd OAI21X1_49/C vdd NAND3X1
XAND2X2_16 INVX1_1/A INVX1_2/A gnd AND2X2_16/Y vdd AND2X2
XNAND3X1_19 INVX1_1/A INVX4_3/A INVX1_32/Y gnd NOR2X1_51/B vdd NAND3X1
XINVX1_32 INVX1_2/A gnd INVX1_32/Y vdd INVX1
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XBUFX2_73 BUFX2_75/A gnd BUFX2_73/Y vdd BUFX2
XBUFX4_8 clk gnd BUFX4_8/Y vdd BUFX4
XBUFX2_64 BUFX2_75/A gnd BUFX2_64/Y vdd BUFX2
XBUFX2_75 BUFX2_75/A gnd BUFX2_75/Y vdd BUFX2
XNOR2X1_29 INVX1_17/Y BUFX4_17/Y gnd NOR2X1_29/Y vdd NOR2X1
XDFFPOSX1_14 BUFX2_29/A BUFX4_8/Y NOR2X1_29/Y gnd vdd DFFPOSX1
XFILL_6_1 gnd vdd FILL
XNAND2X1_9 INVX2_3/A RDATA<2> gnd NAND2X1_9/Y vdd NAND2X1
XBUFX2_22 BUFX2_22/A gnd OUTPD<5> vdd BUFX2
XNAND2X1_12 INVX2_3/A RDATA<3> gnd OAI21X1_8/C vdd NAND2X1
XBUFX2_55 INVX1_6/A gnd WDATA<3> vdd BUFX2
XINVX1_12 INPD<7> gnd INVX1_12/Y vdd INVX1
XAOI21X1_6 INVX2_4/A INVX1_12/Y NOR2X1_2/Y gnd AOI21X1_6/Y vdd AOI21X1
XAOI21X1_1 INVX2_4/A INVX1_7/Y NOR2X1_2/Y gnd OAI21X1_9/C vdd AOI21X1
XNAND2X1_15 INVX2_3/A RDATA<4> gnd OAI21X1_12/C vdd NAND2X1
XOAI21X1_12 INVX2_6/Y INVX2_3/A OAI21X1_12/C gnd OAI21X1_13/A vdd OAI21X1
XOAI21X1_13 OAI21X1_13/A INVX2_4/A AOI21X1_2/Y gnd OAI21X1_14/C vdd OAI21X1
XOAI21X1_14 AND2X2_5/Y OAI21X1_11/Y OAI21X1_14/C gnd OAI21X1_14/Y vdd OAI21X1
XAND2X2_5 AND2X2_5/A INVX2_6/Y gnd AND2X2_5/Y vdd AND2X2
XOAI21X1_11 AND2X2_5/A INVX2_6/Y NOR2X1_2/Y gnd OAI21X1_11/Y vdd OAI21X1
XBUFX4_14 BUFX4_16/A gnd BUFX4_14/Y vdd BUFX4
XNOR2X1_10 NOR2X1_10/A NOR2X1_10/B gnd INVX4_4/A vdd NOR2X1
XDFFPOSX1_22 INVX2_6/A BUFX4_7/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XFILL_5_1_1 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XAOI22X1_2 NOR3X1_1/Y NOR2X1_16/Y AOI22X1_2/C INVX1_8/Y gnd AND2X2_5/A vdd AOI22X1
XNOR2X1_16 INVX1_6/A INVX1_8/Y gnd NOR2X1_16/Y vdd NOR2X1
XINVX1_8 OR2X2_1/B gnd INVX1_8/Y vdd INVX1
XNAND2X1_10 OR2X2_1/B NOR3X1_1/Y gnd OAI21X1_6/C vdd NAND2X1
XOAI21X1_6 OAI21X1_6/A OR2X2_1/B OAI21X1_6/C gnd AND2X2_4/A vdd OAI21X1
XBUFX4_17 BUFX4_16/A gnd BUFX4_17/Y vdd BUFX4
XNOR2X1_2 INVX1_1/A NOR2X1_4/B gnd NOR2X1_2/Y vdd NOR2X1
XNOR2X1_4 NOR2X1_4/A NOR2X1_4/B gnd INVX2_3/A vdd NOR2X1
XNAND2X1_3 OR2X2_1/B INVX1_1/A gnd NOR2X1_4/A vdd NAND2X1
XBUFX4_3 BUFX4_1/A gnd OR2X2_1/B vdd BUFX4
XNAND2X1_2 INVX4_3/A INVX1_2/Y gnd NOR2X1_4/B vdd NAND2X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XNOR2X1_3 INVX4_3/A INVX1_1/A gnd AND2X2_1/A vdd NOR2X1
XAND2X2_1 AND2X2_1/A INVX1_2/Y gnd INVX2_8/A vdd AND2X2
XBUFX4_1 BUFX4_1/A gnd BUFX4_1/Y vdd BUFX4
XXNOR2X1_5 XNOR2X1_5/A BUFX2_5/A gnd XNOR2X1_5/Y vdd XNOR2X1
XFILL_5_0_1 gnd vdd FILL
XFILL_5_0_0 gnd vdd FILL
XXNOR2X1_6 XNOR2X1_6/A BUFX2_6/A gnd XNOR2X1_6/Y vdd XNOR2X1
XNAND2X1_22 INVX2_8/A NAND2X1_22/B gnd XNOR2X1_5/A vdd NAND2X1
XBUFX4_20 BUFX4_22/A gnd BUFX2_75/A vdd BUFX4
XBUFX2_69 BUFX2_75/A gnd BUFX2_69/Y vdd BUFX2
XDFFPOSX1_43 BUFX4_1/A BUFX4_8/Y NAND3X1_20/Y gnd vdd DFFPOSX1
XXOR2X1_3 BUFX2_1/A INVX2_8/A gnd XOR2X1_3/Y vdd XOR2X1
XDFFPOSX1_28 BUFX2_1/A BUFX4_8/Y XOR2X1_3/Y gnd vdd DFFPOSX1
XBUFX2_63 BUFX2_75/A gnd BUFX2_63/Y vdd BUFX2
XINVX1_17 BUFX2_29/A gnd INVX1_17/Y vdd INVX1
XBUFX2_35 BUFX2_75/A gnd PCDELTA<1> vdd BUFX2
XBUFX2_29 BUFX2_29/A gnd OUTPD<12> vdd BUFX2
XFILL_7_1 gnd vdd FILL
XBUFX2_47 BUFX2_44/A gnd PCDELTA<13> vdd BUFX2
XINVX1_7 INPD<3> gnd INVX1_7/Y vdd INVX1
XNAND2X1_19 INVX2_3/A RDATA<7> gnd OAI21X1_28/C vdd NAND2X1
XINVX1_9 INPD<4> gnd INVX1_9/Y vdd INVX1
XOAI21X1_28 INVX2_2/Y INVX2_3/A OAI21X1_28/C gnd OAI21X1_29/A vdd OAI21X1
XOAI21X1_29 OAI21X1_29/A INVX2_4/A AOI21X1_6/Y gnd OAI21X1_30/C vdd OAI21X1
XAOI21X1_2 INVX2_4/A INVX1_9/Y NOR2X1_2/Y gnd AOI21X1_2/Y vdd AOI21X1
XOAI21X1_30 OAI21X1_27/Y AOI21X1_5/Y OAI21X1_30/C gnd OAI21X1_30/Y vdd OAI21X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XOAI21X1_27 AND2X2_10/Y OAI21X1_26/Y NOR2X1_2/Y gnd OAI21X1_27/Y vdd OAI21X1
XNAND3X1_1 INVX4_1/Y INVX2_1/Y NOR2X1_8/Y gnd NOR2X1_10/A vdd NAND3X1
XNOR2X1_8 INVX1_6/A INVX2_6/A gnd NOR2X1_8/Y vdd NOR2X1
XNAND3X1_3 BUFX4_4/Y NOR2X1_8/Y NOR3X1_1/Y gnd NAND3X1_3/Y vdd NAND3X1
XOAI21X1_26 NOR2X1_10/A NOR2X1_10/B BUFX4_4/Y gnd OAI21X1_26/Y vdd OAI21X1
XNAND3X1_2 INVX2_2/Y INVX4_2/Y NOR2X1_9/Y gnd NOR2X1_10/B vdd NAND3X1
XNAND2X1_18 INVX2_1/A INVX2_6/A gnd NOR3X1_3/C vdd NAND2X1
XAND2X2_8 INVX2_1/A INVX2_6/A gnd AND2X2_8/Y vdd AND2X2
XFILL_6_1_1 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XNOR2X1_15 NOR3X1_3/A NOR3X1_3/B gnd AOI22X1_2/C vdd NOR2X1
XNAND2X1_13 INVX1_5/A INVX2_5/A gnd NOR3X1_3/A vdd NAND2X1
XNAND2X1_14 INVX1_6/A INVX4_1/A gnd NOR3X1_3/B vdd NAND2X1
XAND2X2_2 INVX1_5/A INVX2_5/A gnd AND2X2_2/Y vdd AND2X2
XNOR2X1_9 INVX1_5/A INVX2_5/A gnd NOR2X1_9/Y vdd NOR2X1
XNOR3X1_1 INVX1_5/A INVX2_5/A INVX4_1/A gnd NOR3X1_1/Y vdd NOR3X1
XBUFX4_4 BUFX4_1/A gnd BUFX4_4/Y vdd BUFX4
XXNOR2X1_7 XNOR2X1_7/A BUFX2_7/A gnd XNOR2X1_7/Y vdd XNOR2X1
XBUFX4_2 BUFX4_1/A gnd BUFX4_2/Y vdd BUFX4
XNAND2X1_25 OAI21X1_36/Y NAND2X1_25/B gnd XNOR2X1_7/A vdd NAND2X1
XOAI21X1_36 NOR3X1_5/C BUFX2_6/A BUFX4_2/Y gnd OAI21X1_36/Y vdd OAI21X1
XNOR3X1_5 BUFX2_6/A BUFX2_7/A NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XFILL_6_0_1 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XAOI21X1_16 BUFX4_2/Y NOR3X1_5/C INVX2_8/Y gnd NAND2X1_23/B vdd AOI21X1
XNAND2X1_23 OAI21X1_35/Y NAND2X1_23/B gnd XNOR2X1_6/A vdd NAND2X1
XNAND2X1_24 BUFX2_5/A BUFX2_6/A gnd OR2X2_3/A vdd NAND2X1
XINVX1_22 BUFX2_5/A gnd INVX1_22/Y vdd INVX1
XOAI21X1_35 NOR2X1_36/A INVX1_22/Y INVX8_1/Y gnd OAI21X1_35/Y vdd OAI21X1
XNAND3X1_11 INVX2_7/Y INVX1_22/Y NOR3X1_4/Y gnd NOR3X1_5/C vdd NAND3X1
XOAI21X1_34 NOR2X1_36/A OR2X2_2/B NAND3X1_10/Y gnd NAND2X1_22/B vdd OAI21X1
XNAND3X1_10 OR2X2_2/B INVX2_7/Y NOR3X1_4/Y gnd NAND3X1_10/Y vdd NAND3X1
XOAI21X1_33 NOR3X1_4/Y INVX8_1/Y INVX2_8/A gnd AOI21X1_15/C vdd OAI21X1
XAOI21X1_15 INVX8_1/Y AOI21X1_15/B AOI21X1_15/C gnd XNOR2X1_4/A vdd AOI21X1
XXNOR2X1_4 XNOR2X1_4/A INVX2_7/Y gnd XNOR2X1_4/Y vdd XNOR2X1
XINVX2_7 BUFX2_4/A gnd INVX2_7/Y vdd INVX2
XDFFPOSX1_31 BUFX2_4/A BUFX4_8/Y XNOR2X1_4/Y gnd vdd DFFPOSX1
XBUFX2_4 BUFX2_4/A gnd DP<3> vdd BUFX2
XFILL_8_3 gnd vdd FILL
XFILL_8_2 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XBUFX2_56 INVX2_6/A gnd WDATA<4> vdd BUFX2
XAOI21X1_3 INVX2_4/A INVX1_10/Y NOR2X1_2/Y gnd AOI21X1_3/Y vdd AOI21X1
XOAI21X1_18 OAI21X1_17/Y INVX2_4/A AOI21X1_3/Y gnd OAI21X1_19/C vdd OAI21X1
XOAI21X1_17 INVX2_1/Y INVX2_3/A NAND2X1_16/Y gnd OAI21X1_17/Y vdd OAI21X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XOAI21X1_19 AND2X2_7/Y OAI21X1_16/Y OAI21X1_19/C gnd OAI21X1_19/Y vdd OAI21X1
XAND2X2_7 AND2X2_7/A INVX2_1/A gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_16 AND2X2_7/A INVX2_1/A NOR2X1_2/Y gnd OAI21X1_16/Y vdd OAI21X1
XAND2X2_10 NAND3X1_8/Y INVX2_2/A gnd AND2X2_10/Y vdd AND2X2
XAOI21X1_5 AOI21X1_5/A AOI21X1_5/B BUFX4_4/Y gnd AOI21X1_5/Y vdd AOI21X1
XOAI21X1_15 NAND3X1_4/Y BUFX4_4/Y NAND3X1_3/Y gnd AND2X2_7/A vdd OAI21X1
XOAI21X1_25 NAND3X1_6/Y INVX4_2/Y INVX2_2/Y gnd AOI21X1_5/B vdd OAI21X1
XNAND3X1_8 INVX4_2/Y NOR3X1_1/Y NOR3X1_2/Y gnd NAND3X1_8/Y vdd NAND3X1
XNOR3X1_2 INVX1_6/A INVX2_1/A INVX2_6/A gnd NOR3X1_2/Y vdd NOR3X1
XFILL_7_1_1 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XNAND3X1_5 BUFX4_2/Y NOR3X1_1/Y NOR3X1_2/Y gnd NAND3X1_5/Y vdd NAND3X1
XMUX2X1_4 NOR2X1_9/Y AND2X2_2/Y BUFX4_4/Y gnd MUX2X1_4/Y vdd MUX2X1
XNAND3X1_4 INVX2_6/A AND2X2_2/Y AND2X2_6/Y gnd NAND3X1_4/Y vdd NAND3X1
XNAND3X1_6 AND2X2_2/Y AND2X2_6/Y AND2X2_8/Y gnd NAND3X1_6/Y vdd NAND3X1
XAND2X2_6 INVX1_6/A INVX4_1/A gnd AND2X2_6/Y vdd AND2X2
XNAND2X1_11 INVX4_1/A AND2X2_2/Y gnd OAI21X1_6/A vdd NAND2X1
XNOR2X1_14 NOR2X1_9/Y AND2X2_2/Y gnd XNOR2X1_1/A vdd NOR2X1
XXNOR2X1_1 XNOR2X1_1/A BUFX4_4/Y gnd MUX2X1_2/A vdd XNOR2X1
XDFFPOSX1_34 BUFX2_7/A BUFX4_12/Y XNOR2X1_7/Y gnd vdd DFFPOSX1
XINVX8_1 BUFX4_2/Y gnd INVX8_1/Y vdd INVX8
XAOI21X1_17 INVX8_1/Y INVX1_23/Y INVX2_8/Y gnd NAND2X1_25/B vdd AOI21X1
XAOI21X1_18 INVX8_1/Y NAND2X1_26/Y INVX2_8/Y gnd AOI21X1_18/Y vdd AOI21X1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XFILL_7_0_1 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XNAND2X1_26 BUFX2_7/A INVX1_23/A gnd NAND2X1_26/Y vdd NAND2X1
XNOR2X1_38 INVX2_8/Y NOR2X1_37/Y gnd NOR2X1_38/Y vdd NOR2X1
XNAND2X1_27 BUFX2_7/A BUFX2_8/A gnd OR2X2_3/B vdd NAND2X1
XNOR2X1_35 OR2X2_3/A NOR2X1_36/A gnd INVX1_23/A vdd NOR2X1
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XNOR2X1_36 NOR2X1_36/A OR2X2_3/Y gnd NOR2X1_37/B vdd NOR2X1
XNOR2X1_37 OR2X2_2/B NOR2X1_37/B gnd NOR2X1_37/Y vdd NOR2X1
XBUFX4_6 BUFX4_1/A gnd OR2X2_2/B vdd BUFX4
XNAND2X1_21 AND2X2_12/Y OR2X2_2/A gnd NOR2X1_36/A vdd NAND2X1
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XNAND3X1_9 INVX2_8/A NAND3X1_9/B OR2X2_2/Y gnd XNOR2X1_3/A vdd NAND3X1
XNAND2X1_20 BUFX2_3/A OR2X2_2/A gnd AOI21X1_15/B vdd NAND2X1
XAND2X2_11 BUFX2_1/A BUFX2_2/A gnd OR2X2_2/A vdd AND2X2
XAND2X2_12 BUFX2_3/A BUFX2_4/A gnd AND2X2_12/Y vdd AND2X2
XNOR3X1_4 BUFX2_1/A BUFX2_2/A BUFX2_3/A gnd NOR3X1_4/Y vdd NOR3X1
XBUFX2_1 BUFX2_1/A gnd DP<0> vdd BUFX2
XFILL_9_1 gnd vdd FILL
XBUFX2_59 INVX2_2/A gnd WDATA<7> vdd BUFX2
XBUFX4_18 BUFX4_22/A gnd BUFX2_44/A vdd BUFX4
XDFFPOSX1_25 INVX2_2/A BUFX4_11/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_23 INVX2_1/A BUFX4_11/Y OAI21X1_19/Y gnd vdd DFFPOSX1
XINVX4_2 INVX4_2/A gnd INVX4_2/Y vdd INVX4
XNAND3X1_7 INVX2_2/A INVX4_2/A NOR3X1_3/Y gnd AOI21X1_5/A vdd NAND3X1
XOAI22X1_1 NOR2X1_2/Y MUX2X1_3/Y AND2X2_3/Y OAI21X1_5/Y gnd OAI22X1_1/Y vdd OAI22X1
XAND2X2_3 MUX2X1_4/Y INVX4_1/Y gnd AND2X2_3/Y vdd AND2X2
XOAI21X1_5 MUX2X1_4/Y INVX4_1/Y NOR2X1_2/Y gnd OAI21X1_5/Y vdd OAI21X1
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XBUFX4_11 clk gnd BUFX4_11/Y vdd BUFX4
XFILL_8_1_1 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XOAI21X1_20 NAND3X1_6/Y BUFX4_2/Y NAND3X1_5/Y gnd AND2X2_9/A vdd OAI21X1
XBUFX4_12 clk gnd BUFX4_12/Y vdd BUFX4
XBUFX2_74 BUFX2_70/A gnd BUFX2_74/Y vdd BUFX2
XBUFX4_19 BUFX4_22/A gnd BUFX2_70/A vdd BUFX4
XDFFPOSX1_35 BUFX2_8/A BUFX4_12/Y XNOR2X1_8/Y gnd vdd DFFPOSX1
XXNOR2X1_8 XNOR2X1_8/A BUFX2_8/A gnd XNOR2X1_8/Y vdd XNOR2X1
XBUFX4_5 BUFX4_1/A gnd BUFX4_5/Y vdd BUFX4
XOAI21X1_37 INVX8_1/Y NOR3X1_5/Y AOI21X1_18/Y gnd XNOR2X1_8/A vdd OAI21X1
XINVX1_24 BUFX2_8/A gnd INVX1_24/Y vdd INVX1
XAND2X2_13 NOR3X1_5/Y INVX1_24/Y gnd AND2X2_13/Y vdd AND2X2
XNAND3X1_12 INVX1_24/Y INVX1_25/Y NOR3X1_5/Y gnd NOR3X1_6/C vdd NAND3X1
XINVX1_25 BUFX2_9/A gnd INVX1_25/Y vdd INVX1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XOAI21X1_39 BUFX4_5/Y BUFX2_9/A NOR2X1_38/Y gnd AOI21X1_19/C vdd OAI21X1
XOAI21X1_38 AND2X2_13/Y INVX8_1/Y NOR2X1_38/Y gnd XNOR2X1_9/A vdd OAI21X1
XFILL_8_0_1 gnd vdd FILL
XFILL_8_0_0 gnd vdd FILL
XNAND3X1_13 BUFX2_9/A XOR2X1_4/B NOR2X1_37/B gnd NOR3X1_7/C vdd NAND3X1
XDFFPOSX1_37 XOR2X1_4/B BUFX4_9/Y XOR2X1_4/Y gnd vdd DFFPOSX1
XXNOR2X1_9 XNOR2X1_9/A BUFX2_9/A gnd XNOR2X1_9/Y vdd XNOR2X1
XNOR2X1_33 OR2X2_2/B INVX1_21/Y gnd NOR2X1_33/Y vdd NOR2X1
XINVX1_21 BUFX2_1/A gnd INVX1_21/Y vdd INVX1
XBUFX4_9 clk gnd BUFX4_9/Y vdd BUFX4
XOAI21X1_32 BUFX2_1/A BUFX2_2/A OR2X2_2/B gnd NAND3X1_9/B vdd OAI21X1
XXNOR2X1_3 XNOR2X1_3/A BUFX2_3/A gnd XNOR2X1_3/Y vdd XNOR2X1
XDFFPOSX1_36 BUFX2_9/A BUFX4_9/Y XNOR2X1_9/Y gnd vdd DFFPOSX1
XBUFX2_9 BUFX2_9/A gnd DP<8> vdd BUFX2
XFILL_10_2 gnd vdd FILL
XFILL_10_1 gnd vdd FILL
XBUFX2_44 BUFX2_44/A gnd PCDELTA<10> vdd BUFX2
XINVX1_11 INPD<6> gnd INVX1_11/Y vdd INVX1
XBUFX2_58 INVX4_2/A gnd WDATA<6> vdd BUFX2
XAOI21X1_4 INVX2_4/A INVX1_11/Y NOR2X1_2/Y gnd AOI21X1_4/Y vdd AOI21X1
XDFFPOSX1_24 INVX4_2/A BUFX4_11/Y OAI21X1_24/Y gnd vdd DFFPOSX1
XOAI21X1_23 OAI21X1_22/Y INVX2_4/A AOI21X1_4/Y gnd OAI21X1_24/C vdd OAI21X1
XOAI21X1_24 AND2X2_9/Y OAI21X1_21/Y OAI21X1_24/C gnd OAI21X1_24/Y vdd OAI21X1
XAND2X2_9 AND2X2_9/A INVX4_2/A gnd AND2X2_9/Y vdd AND2X2
XOAI21X1_21 AND2X2_9/A INVX4_2/A NOR2X1_2/Y gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_22 INVX4_2/Y INVX2_3/A OAI21X1_22/C gnd OAI21X1_22/Y vdd OAI21X1
XDFFPOSX1_20 INVX4_1/A BUFX4_11/Y OAI22X1_1/Y gnd vdd DFFPOSX1
XBUFX2_54 INVX4_1/A gnd WDATA<2> vdd BUFX2
XFILL_9_1_1 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XNOR2X1_13 NOR2X1_2/Y INVX2_4/Y gnd XOR2X1_2/A vdd NOR2X1
XBUFX2_71 BUFX2_70/A gnd BUFX2_71/Y vdd BUFX2
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B NOR2X1_2/Y gnd MUX2X1_2/Y vdd MUX2X1
XBUFX2_70 BUFX2_70/A gnd BUFX2_70/Y vdd BUFX2
XBUFX2_61 BUFX4_2/Y gnd BUFX2_61/Y vdd BUFX2
XDFFPOSX1_16 INVX1_19/A BUFX4_12/Y NOR2X1_31/Y gnd vdd DFFPOSX1
XNOR2X1_31 INVX1_19/Y BUFX4_17/Y gnd NOR2X1_31/Y vdd NOR2X1
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XOAI21X1_44 BUFX4_2/Y INVX1_28/A OAI21X1_44/C gnd AOI21X1_22/C vdd OAI21X1
XAOI21X1_22 BUFX4_5/Y INVX1_28/A AOI21X1_22/C gnd NAND3X1_14/C vdd AOI21X1
XBUFX2_8 BUFX2_8/A gnd DP<7> vdd BUFX2
XNAND3X1_14 INVX2_8/A NAND3X1_14/B NAND3X1_14/C gnd INVX1_29/A vdd NAND3X1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XAOI21X1_19 BUFX4_5/Y NOR3X1_6/C AOI21X1_19/C gnd XOR2X1_4/A vdd AOI21X1
XAOI21X1_20 INVX8_1/Y NOR3X1_7/C INVX2_8/Y gnd OAI21X1_40/C vdd AOI21X1
XFILL_9_0_1 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XOAI21X1_40 NOR2X1_39/Y INVX8_1/Y OAI21X1_40/C gnd XNOR2X1_10/A vdd OAI21X1
XNOR2X1_39 XOR2X1_4/B NOR3X1_6/C gnd NOR2X1_39/Y vdd NOR2X1
XXOR2X1_4 XOR2X1_4/A XOR2X1_4/B gnd XOR2X1_4/Y vdd XOR2X1
XNOR2X1_34 BUFX2_1/A INVX8_1/Y gnd NOR2X1_34/Y vdd NOR2X1
XOAI21X1_31 NOR2X1_33/Y NOR2X1_34/Y INVX2_8/A gnd XNOR2X1_2/A vdd OAI21X1
XXNOR2X1_2 XNOR2X1_2/A BUFX2_2/A gnd XNOR2X1_2/Y vdd XNOR2X1
XDFFPOSX1_29 BUFX2_2/A BUFX4_9/Y XNOR2X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_30 BUFX2_3/A BUFX4_9/Y XNOR2X1_3/Y gnd vdd DFFPOSX1
XBUFX2_3 BUFX2_3/A gnd DP<2> vdd BUFX2
XBUFX2_2 BUFX2_2/A gnd DP<1> vdd BUFX2
XDFFPOSX1_13 INVX1_16/A BUFX4_11/Y NOR2X1_28/Y gnd vdd DFFPOSX1
XNOR2X1_28 INVX1_16/Y BUFX4_14/Y gnd NOR2X1_28/Y vdd NOR2X1
XNOR2X1_19 BUFX2_19/A BUFX4_14/Y gnd AOI21X1_9/C vdd NOR2X1
XAOI21X1_9 INVX4_1/Y BUFX4_14/Y AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XOAI21X1_4 INVX4_1/Y INVX2_3/A NAND2X1_9/Y gnd MUX2X1_3/A vdd OAI21X1
XNOR2X1_18 BUFX2_18/A BUFX4_14/Y gnd AOI21X1_8/C vdd NOR2X1
XAOI21X1_8 INVX1_5/Y BUFX4_14/Y AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XMUX2X1_3 MUX2X1_3/A INPD<2> INVX2_4/Y gnd MUX2X1_3/Y vdd MUX2X1
XOAI21X1_3 INVX1_5/Y INVX2_3/A OAI21X1_3/C gnd MUX2X1_1/A vdd OAI21X1
XMUX2X1_1 MUX2X1_1/A INPD<1> INVX2_4/Y gnd MUX2X1_2/B vdd MUX2X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XDFFPOSX1_26 XOR2X1_2/B BUFX4_12/Y XOR2X1_2/Y gnd vdd DFFPOSX1
XFILL_10_1_1 gnd vdd FILL
XFILL_10_1_0 gnd vdd FILL
XDFFPOSX1_19 INVX1_5/A BUFX4_12/Y MUX2X1_2/Y gnd vdd DFFPOSX1
XBUFX2_31 INVX1_19/A gnd OUTPD<14> vdd BUFX2
XDFFPOSX1_41 INVX1_28/A BUFX4_12/Y XNOR2X1_13/Y gnd vdd DFFPOSX1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XXNOR2X1_13 NOR3X1_8/Y INVX1_28/Y gnd XNOR2X1_13/Y vdd XNOR2X1
XNAND2X1_29 BUFX4_5/Y INVX2_9/A gnd OAI21X1_44/C vdd NAND2X1
XNAND2X1_30 OAI21X1_44/C NAND3X1_14/B gnd NOR3X1_8/B vdd NAND2X1
XOAI21X1_43 NOR3X1_7/Y BUFX4_5/Y INVX2_8/A gnd NOR3X1_8/A vdd OAI21X1
XOAI21X1_45 NOR3X1_7/Y BUFX4_5/Y INVX1_29/Y gnd NOR2X1_41/A vdd OAI21X1
XNOR3X1_7 INVX1_26/Y NOR3X1_7/B NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XFILL_10_0_1 gnd vdd FILL
XFILL_10_0_0 gnd vdd FILL
XOAI21X1_41 NOR3X1_7/C INVX1_26/Y INVX8_1/Y gnd AND2X2_14/A vdd OAI21X1
XAND2X2_14 AND2X2_14/A INVX2_8/A gnd AND2X2_14/Y vdd AND2X2
XINVX1_26 BUFX2_11/A gnd INVX1_26/Y vdd INVX1
XNOR3X1_6 XOR2X1_4/B BUFX2_11/A NOR3X1_6/C gnd NOR3X1_6/Y vdd NOR3X1
XXNOR2X1_10 XNOR2X1_10/A BUFX2_11/A gnd XNOR2X1_10/Y vdd XNOR2X1
XDFFPOSX1_38 BUFX2_11/A BUFX4_9/Y XNOR2X1_10/Y gnd vdd DFFPOSX1
XBUFX2_11 BUFX2_11/A gnd DP<10> vdd BUFX2
XNOR2X1_27 INVX1_15/Y BUFX4_17/Y gnd NOR2X1_27/Y vdd NOR2X1
XINVX1_15 BUFX2_27/A gnd INVX1_15/Y vdd INVX1
XDFFPOSX1_12 BUFX2_27/A BUFX4_9/Y NOR2X1_27/Y gnd vdd DFFPOSX1
XBUFX2_27 BUFX2_27/A gnd OUTPD<10> vdd BUFX2
XFILL_12_1 gnd vdd FILL
XBUFX2_48 BUFX2_44/A gnd PCDELTA<14> vdd BUFX2
XBUFX2_36 BUFX2_44/A gnd PCDELTA<2> vdd BUFX2
XBUFX2_45 BUFX2_44/A gnd PCDELTA<11> vdd BUFX2
XBUFX2_65 BUFX2_44/A gnd BUFX2_65/Y vdd BUFX2
XBUFX2_28 INVX1_16/A gnd OUTPD<11> vdd BUFX2
XDFFPOSX1_4 BUFX2_19/A BUFX4_11/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XBUFX2_19 BUFX2_19/A gnd OUTPD<2> vdd BUFX2
XBUFX2_18 BUFX2_18/A gnd OUTPD<1> vdd BUFX2
XDFFPOSX1_3 BUFX2_18/A BUFX4_11/Y AOI21X1_8/Y gnd vdd DFFPOSX1
XNAND2X1_17 INVX2_3/A RDATA<6> gnd OAI21X1_22/C vdd NAND2X1
XNAND2X1_8 INVX2_3/A RDATA<1> gnd OAI21X1_3/C vdd NAND2X1
XBUFX2_57 INVX2_1/A gnd WDATA<5> vdd BUFX2
XBUFX2_16 XOR2X1_2/B gnd IR vdd BUFX2
XFILL_11_1_1 gnd vdd FILL
XFILL_11_1_0 gnd vdd FILL
XXOR2X1_2 XOR2X1_2/A XOR2X1_2/B gnd XOR2X1_2/Y vdd XOR2X1
XBUFX2_53 INVX1_5/A gnd WDATA<1> vdd BUFX2
XBUFX2_39 BUFX2_70/A gnd PCDELTA<5> vdd BUFX2
XBUFX2_37 BUFX2_70/A gnd PCDELTA<3> vdd BUFX2
XBUFX2_49 BUFX2_70/A gnd PCDELTA<15> vdd BUFX2
XBUFX2_7 BUFX2_7/A gnd DP<6> vdd BUFX2
XBUFX2_13 INVX2_9/A gnd DP<12> vdd BUFX2
XDFFPOSX1_40 INVX2_9/A BUFX4_12/Y XNOR2X1_12/Y gnd vdd DFFPOSX1
XBUFX2_14 INVX1_28/A gnd DP<13> vdd BUFX2
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XNAND2X1_28 INVX8_1/Y INVX2_9/Y gnd NAND3X1_14/B vdd NAND2X1
XXNOR2X1_12 NOR2X1_40/Y INVX2_9/Y gnd XNOR2X1_12/Y vdd XNOR2X1
XNOR2X1_40 NOR3X1_8/A NOR3X1_8/C gnd NOR2X1_40/Y vdd NOR2X1
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd NOR3X1_8/Y vdd NOR3X1
XFILL_11_0_1 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XBUFX2_10 XOR2X1_4/B gnd DP<9> vdd BUFX2
XNOR2X1_41 NOR2X1_41/A NOR3X1_8/C gnd XOR2X1_5/A vdd NOR2X1
XAOI21X1_21 NOR3X1_7/B NOR3X1_6/Y INVX8_1/Y gnd NOR3X1_8/C vdd AOI21X1
XOAI21X1_42 INVX8_1/Y NOR3X1_6/Y AND2X2_14/Y gnd XNOR2X1_11/A vdd OAI21X1
XXOR2X1_5 XOR2X1_5/A BUFX2_15/A gnd XOR2X1_5/Y vdd XOR2X1
XDFFPOSX1_42 BUFX2_15/A BUFX4_9/Y XOR2X1_5/Y gnd vdd DFFPOSX1
XBUFX2_15 BUFX2_15/A gnd DP<14> vdd BUFX2
XINVX1_27 BUFX2_12/A gnd NOR3X1_7/B vdd INVX1
XXNOR2X1_11 XNOR2X1_11/A BUFX2_12/A gnd XNOR2X1_11/Y vdd XNOR2X1
XBUFX2_12 BUFX2_12/A gnd DP<11> vdd BUFX2
XDFFPOSX1_39 BUFX2_12/A BUFX4_9/Y XNOR2X1_11/Y gnd vdd DFFPOSX1
.ends

