VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO BFCPU
   FOREIGN BFCPU ;
   ORIGIN 2.6000 3.0000 ;
   SIZE 153.9000 BY 126.1000 ;
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 0.2000 120.2000 148.6000 120.8000 ;
	    RECT 1.4000 115.9000 1.8000 120.2000 ;
	    RECT 4.2000 117.9000 4.6000 120.2000 ;
	    RECT 5.8000 117.9000 6.2000 120.2000 ;
	    RECT 8.6000 116.0000 9.0000 120.2000 ;
	    RECT 11.0000 116.5000 11.4000 120.2000 ;
	    RECT 13.4000 116.6000 13.9000 120.2000 ;
	    RECT 16.5000 119.9000 16.9000 120.2000 ;
	    RECT 16.5000 116.6000 17.0000 119.9000 ;
	    RECT 18.2000 117.9000 18.6000 120.2000 ;
	    RECT 20.6000 116.5000 21.0000 120.2000 ;
	    RECT 23.0000 115.9000 23.4000 120.2000 ;
	    RECT 25.8000 117.9000 26.2000 120.2000 ;
	    RECT 27.4000 117.9000 27.8000 120.2000 ;
	    RECT 30.2000 116.0000 30.6000 120.2000 ;
	    RECT 32.6000 116.6000 33.1000 120.2000 ;
	    RECT 35.7000 119.9000 36.1000 120.2000 ;
	    RECT 35.7000 116.6000 36.2000 119.9000 ;
	    RECT 37.4000 115.9000 37.8000 120.2000 ;
	    RECT 39.5000 117.9000 39.9000 120.2000 ;
	    RECT 41.4000 116.5000 41.8000 120.2000 ;
	    RECT 45.4000 115.9000 45.8000 120.2000 ;
	    RECT 47.0000 116.5000 47.4000 120.2000 ;
	    RECT 55.0000 116.9000 55.4000 120.2000 ;
	    RECT 58.2000 115.9000 58.6000 120.2000 ;
	    RECT 59.9000 119.9000 60.3000 120.2000 ;
	    RECT 59.8000 116.6000 60.3000 119.9000 ;
	    RECT 62.9000 116.6000 63.4000 120.2000 ;
	    RECT 64.6000 117.9000 65.0000 120.2000 ;
	    RECT 66.2000 117.9000 66.6000 120.2000 ;
	    RECT 67.8000 115.9000 68.2000 120.2000 ;
	    RECT 69.4000 116.5000 69.8000 120.2000 ;
	    RECT 71.8000 116.0000 72.2000 120.2000 ;
	    RECT 74.6000 117.9000 75.0000 120.2000 ;
	    RECT 76.2000 117.9000 76.6000 120.2000 ;
	    RECT 79.0000 115.9000 79.4000 120.2000 ;
	    RECT 81.4000 116.5000 81.8000 120.2000 ;
	    RECT 83.8000 116.5000 84.2000 120.2000 ;
	    RECT 86.2000 116.5000 86.6000 120.2000 ;
	    RECT 88.6000 116.5000 89.0000 120.2000 ;
	    RECT 91.0000 116.5000 91.4000 120.2000 ;
	    RECT 93.4000 116.5000 93.8000 120.2000 ;
	    RECT 95.9000 119.9000 96.3000 120.2000 ;
	    RECT 95.8000 116.6000 96.3000 119.9000 ;
	    RECT 98.9000 116.6000 99.4000 120.2000 ;
	    RECT 103.0000 116.5000 103.4000 120.2000 ;
	    RECT 105.4000 116.5000 105.8000 120.2000 ;
	    RECT 107.0000 117.9000 107.4000 120.2000 ;
	    RECT 108.6000 117.9000 109.0000 120.2000 ;
	    RECT 109.4000 117.9000 109.8000 120.2000 ;
	    RECT 111.0000 117.9000 111.4000 120.2000 ;
	    RECT 112.6000 116.0000 113.0000 120.2000 ;
	    RECT 115.4000 117.9000 115.8000 120.2000 ;
	    RECT 117.0000 117.9000 117.4000 120.2000 ;
	    RECT 119.8000 115.9000 120.2000 120.2000 ;
	    RECT 122.2000 116.5000 122.6000 120.2000 ;
	    RECT 124.6000 116.5000 125.0000 120.2000 ;
	    RECT 127.0000 115.9000 127.4000 120.2000 ;
	    RECT 129.8000 117.9000 130.2000 120.2000 ;
	    RECT 131.4000 117.9000 131.8000 120.2000 ;
	    RECT 134.2000 116.0000 134.6000 120.2000 ;
	    RECT 136.6000 116.5000 137.0000 120.2000 ;
	    RECT 139.0000 116.5000 139.4000 120.2000 ;
	    RECT 141.4000 116.5000 141.8000 120.2000 ;
	    RECT 143.8000 116.5000 144.2000 120.2000 ;
	    RECT 146.2000 116.5000 146.6000 120.2000 ;
	    RECT 1.4000 100.8000 1.8000 104.5000 ;
	    RECT 3.8000 100.8000 4.2000 105.1000 ;
	    RECT 6.6000 100.8000 7.0000 103.1000 ;
	    RECT 8.2000 100.8000 8.6000 103.1000 ;
	    RECT 11.0000 100.8000 11.4000 105.0000 ;
	    RECT 12.6000 100.8000 13.0000 103.1000 ;
	    RECT 14.2000 100.8000 14.6000 105.1000 ;
	    RECT 17.4000 100.8000 17.8000 104.5000 ;
	    RECT 19.8000 100.8000 20.2000 105.1000 ;
	    RECT 22.6000 100.8000 23.0000 103.1000 ;
	    RECT 24.2000 100.8000 24.6000 103.1000 ;
	    RECT 27.0000 100.8000 27.4000 105.0000 ;
	    RECT 29.4000 100.8000 29.9000 104.4000 ;
	    RECT 32.5000 101.1000 33.0000 104.4000 ;
	    RECT 32.5000 100.8000 32.9000 101.1000 ;
	    RECT 39.0000 100.8000 39.4000 104.1000 ;
	    RECT 40.6000 100.8000 41.0000 103.1000 ;
	    RECT 43.0000 100.8000 43.4000 104.9000 ;
	    RECT 44.6000 100.8000 45.0000 103.1000 ;
	    RECT 45.7000 100.8000 46.1000 103.1000 ;
	    RECT 47.8000 100.8000 48.2000 105.1000 ;
	    RECT 51.0000 100.8000 51.4000 104.1000 ;
	    RECT 56.9000 100.8000 57.3000 103.1000 ;
	    RECT 59.0000 100.8000 59.4000 105.1000 ;
	    RECT 60.1000 100.8000 60.5000 103.1000 ;
	    RECT 62.2000 100.8000 62.6000 105.1000 ;
	    RECT 63.0000 100.8000 63.4000 103.1000 ;
	    RECT 64.6000 100.8000 65.0000 103.1000 ;
	    RECT 65.4000 100.8000 65.8000 103.1000 ;
	    RECT 67.0000 100.8000 67.4000 103.1000 ;
	    RECT 68.6000 101.1000 69.1000 104.4000 ;
	    RECT 68.7000 100.8000 69.1000 101.1000 ;
	    RECT 71.7000 100.8000 72.2000 104.4000 ;
	    RECT 74.2000 100.8000 74.6000 103.1000 ;
	    RECT 75.8000 100.8000 76.2000 105.1000 ;
	    RECT 78.6000 100.8000 79.0000 103.1000 ;
	    RECT 80.2000 100.8000 80.6000 103.1000 ;
	    RECT 83.0000 100.8000 83.4000 105.0000 ;
	    RECT 85.4000 100.8000 85.8000 104.5000 ;
	    RECT 87.8000 100.8000 88.2000 105.0000 ;
	    RECT 90.6000 100.8000 91.0000 103.1000 ;
	    RECT 92.2000 100.8000 92.6000 103.1000 ;
	    RECT 95.0000 100.8000 95.4000 105.1000 ;
	    RECT 99.0000 100.8000 99.4000 105.0000 ;
	    RECT 101.8000 100.8000 102.2000 103.1000 ;
	    RECT 103.4000 100.8000 103.8000 103.1000 ;
	    RECT 106.2000 100.8000 106.6000 105.1000 ;
	    RECT 107.8000 100.8000 108.2000 103.1000 ;
	    RECT 110.2000 100.8000 110.6000 104.9000 ;
	    RECT 112.8000 100.8000 113.2000 105.1000 ;
	    RECT 114.5000 100.8000 114.9000 103.1000 ;
	    RECT 116.6000 100.8000 117.0000 105.1000 ;
	    RECT 118.2000 100.8000 118.6000 104.9000 ;
	    RECT 120.8000 100.8000 121.2000 105.1000 ;
	    RECT 123.0000 100.8000 123.4000 104.5000 ;
	    RECT 125.4000 100.8000 125.8000 105.1000 ;
	    RECT 127.8000 100.8000 128.2000 105.1000 ;
	    RECT 129.9000 100.8000 130.3000 103.1000 ;
	    RECT 131.8000 100.8000 132.2000 104.5000 ;
	    RECT 134.2000 100.8000 134.6000 105.1000 ;
	    RECT 138.2000 100.8000 138.6000 105.1000 ;
	    RECT 139.8000 100.8000 140.2000 105.0000 ;
	    RECT 142.6000 100.8000 143.0000 103.1000 ;
	    RECT 144.2000 100.8000 144.6000 103.1000 ;
	    RECT 147.0000 100.8000 147.4000 105.1000 ;
	    RECT 0.2000 100.2000 148.6000 100.8000 ;
	    RECT 1.4000 96.5000 1.8000 100.2000 ;
	    RECT 3.8000 96.5000 4.2000 100.2000 ;
	    RECT 6.2000 95.9000 6.6000 100.2000 ;
	    RECT 9.0000 97.9000 9.4000 100.2000 ;
	    RECT 10.6000 97.9000 11.0000 100.2000 ;
	    RECT 13.4000 96.0000 13.8000 100.2000 ;
	    RECT 15.8000 95.9000 16.2000 100.2000 ;
	    RECT 18.6000 97.9000 19.0000 100.2000 ;
	    RECT 20.2000 97.9000 20.6000 100.2000 ;
	    RECT 23.0000 96.0000 23.4000 100.2000 ;
	    RECT 25.4000 96.6000 25.9000 100.2000 ;
	    RECT 28.5000 99.9000 28.9000 100.2000 ;
	    RECT 28.5000 96.6000 29.0000 99.9000 ;
	    RECT 30.2000 95.9000 30.6000 100.2000 ;
	    RECT 32.3000 97.9000 32.7000 100.2000 ;
	    RECT 33.4000 95.9000 33.8000 100.2000 ;
	    RECT 36.6000 96.6000 37.1000 100.2000 ;
	    RECT 39.7000 99.9000 40.1000 100.2000 ;
	    RECT 39.7000 96.6000 40.2000 99.9000 ;
	    RECT 43.0000 95.9000 43.4000 100.2000 ;
	    RECT 43.8000 95.9000 44.2000 100.2000 ;
	    RECT 45.9000 97.9000 46.3000 100.2000 ;
	    RECT 50.2000 96.5000 50.6000 100.2000 ;
	    RECT 53.4000 96.5000 53.8000 100.2000 ;
	    RECT 55.8000 97.9000 56.2000 100.2000 ;
	    RECT 56.6000 97.9000 57.0000 100.2000 ;
	    RECT 58.2000 98.1000 58.6000 100.2000 ;
	    RECT 60.6000 96.5000 61.0000 100.2000 ;
	    RECT 63.0000 96.5000 63.4000 100.2000 ;
	    RECT 65.7000 97.9000 66.1000 100.2000 ;
	    RECT 67.8000 95.9000 68.2000 100.2000 ;
	    RECT 68.6000 97.9000 69.0000 100.2000 ;
	    RECT 70.2000 95.9000 70.6000 100.2000 ;
	    RECT 73.4000 96.0000 73.8000 100.2000 ;
	    RECT 76.2000 97.9000 76.6000 100.2000 ;
	    RECT 77.8000 97.9000 78.2000 100.2000 ;
	    RECT 80.6000 95.9000 81.0000 100.2000 ;
	    RECT 83.0000 96.5000 83.4000 100.2000 ;
	    RECT 85.4000 96.5000 85.8000 100.2000 ;
	    RECT 87.6000 95.9000 88.0000 100.2000 ;
	    RECT 90.2000 96.1000 90.6000 100.2000 ;
	    RECT 92.6000 96.5000 93.0000 100.2000 ;
	    RECT 94.2000 95.9000 94.6000 100.2000 ;
	    RECT 97.4000 95.9000 97.8000 100.2000 ;
	    RECT 100.6000 96.5000 101.0000 100.2000 ;
	    RECT 103.0000 95.9000 103.4000 100.2000 ;
	    RECT 105.8000 97.9000 106.2000 100.2000 ;
	    RECT 107.4000 97.9000 107.8000 100.2000 ;
	    RECT 110.2000 96.0000 110.6000 100.2000 ;
	    RECT 112.1000 97.9000 112.5000 100.2000 ;
	    RECT 114.2000 95.9000 114.6000 100.2000 ;
	    RECT 115.3000 97.9000 115.7000 100.2000 ;
	    RECT 117.4000 95.9000 117.8000 100.2000 ;
	    RECT 118.2000 97.9000 118.6000 100.2000 ;
	    RECT 119.8000 96.1000 120.2000 100.2000 ;
	    RECT 121.4000 95.9000 121.8000 100.2000 ;
	    RECT 123.5000 97.9000 123.9000 100.2000 ;
	    RECT 124.6000 95.9000 125.0000 100.2000 ;
	    RECT 126.7000 97.9000 127.1000 100.2000 ;
	    RECT 128.6000 96.0000 129.0000 100.2000 ;
	    RECT 131.4000 97.9000 131.8000 100.2000 ;
	    RECT 133.0000 97.9000 133.4000 100.2000 ;
	    RECT 135.8000 95.9000 136.2000 100.2000 ;
	    RECT 139.0000 96.5000 139.4000 100.2000 ;
	    RECT 141.4000 96.5000 141.8000 100.2000 ;
	    RECT 143.8000 97.9000 144.2000 100.2000 ;
	    RECT 145.4000 96.5000 145.8000 100.2000 ;
	    RECT 1.4000 80.8000 1.8000 84.5000 ;
	    RECT 3.8000 80.8000 4.2000 85.1000 ;
	    RECT 6.6000 80.8000 7.0000 83.1000 ;
	    RECT 8.2000 80.8000 8.6000 83.1000 ;
	    RECT 11.0000 80.8000 11.4000 85.0000 ;
	    RECT 13.4000 80.8000 13.9000 84.4000 ;
	    RECT 16.5000 81.1000 17.0000 84.4000 ;
	    RECT 16.5000 80.8000 16.9000 81.1000 ;
	    RECT 18.2000 80.8000 18.6000 85.1000 ;
	    RECT 20.3000 80.8000 20.7000 83.1000 ;
	    RECT 22.2000 80.8000 22.6000 84.5000 ;
	    RECT 23.8000 80.8000 24.2000 85.1000 ;
	    RECT 24.6000 80.8000 25.0000 83.1000 ;
	    RECT 27.8000 80.8000 28.2000 85.1000 ;
	    RECT 29.4000 80.8000 29.9000 84.4000 ;
	    RECT 32.5000 81.1000 33.0000 84.4000 ;
	    RECT 32.5000 80.8000 32.9000 81.1000 ;
	    RECT 35.0000 80.8000 35.4000 85.0000 ;
	    RECT 37.8000 80.8000 38.2000 83.1000 ;
	    RECT 39.4000 80.8000 39.8000 83.1000 ;
	    RECT 42.2000 80.8000 42.6000 85.1000 ;
	    RECT 44.6000 80.8000 45.0000 82.9000 ;
	    RECT 46.2000 80.8000 46.6000 83.1000 ;
	    RECT 48.9000 80.8000 49.3000 83.1000 ;
	    RECT 51.0000 80.8000 51.4000 85.1000 ;
	    RECT 52.1000 80.8000 52.5000 83.1000 ;
	    RECT 54.2000 80.8000 54.6000 85.1000 ;
	    RECT 55.8000 80.8000 56.2000 85.1000 ;
	    RECT 56.6000 80.8000 57.0000 83.1000 ;
	    RECT 59.0000 80.8000 59.4000 82.9000 ;
	    RECT 60.6000 80.8000 61.0000 83.1000 ;
	    RECT 62.2000 80.8000 62.6000 84.9000 ;
	    RECT 63.8000 80.8000 64.2000 83.1000 ;
	    RECT 65.4000 80.8000 65.8000 83.1000 ;
	    RECT 66.2000 80.8000 66.6000 85.1000 ;
	    RECT 68.3000 80.8000 68.7000 83.1000 ;
	    RECT 69.4000 80.8000 69.8000 85.1000 ;
	    RECT 71.0000 80.8000 71.4000 84.5000 ;
	    RECT 73.4000 81.1000 73.9000 84.4000 ;
	    RECT 73.5000 80.8000 73.9000 81.1000 ;
	    RECT 76.5000 80.8000 77.0000 84.4000 ;
	    RECT 79.0000 80.8000 79.4000 85.1000 ;
	    RECT 81.8000 80.8000 82.2000 83.1000 ;
	    RECT 83.4000 80.8000 83.8000 83.1000 ;
	    RECT 86.2000 80.8000 86.6000 85.0000 ;
	    RECT 88.6000 80.8000 89.0000 84.5000 ;
	    RECT 90.2000 80.8000 90.6000 85.1000 ;
	    RECT 91.8000 80.8000 92.2000 84.5000 ;
	    RECT 94.2000 80.8000 94.6000 84.5000 ;
	    RECT 95.8000 80.8000 96.2000 85.1000 ;
	    RECT 96.9000 80.8000 97.3000 83.1000 ;
	    RECT 99.0000 80.8000 99.4000 85.1000 ;
	    RECT 102.2000 80.8000 102.6000 84.5000 ;
	    RECT 103.8000 80.8000 104.2000 85.1000 ;
	    RECT 104.6000 80.8000 105.0000 85.1000 ;
	    RECT 106.2000 80.8000 106.6000 85.1000 ;
	    RECT 107.0000 80.8000 107.4000 85.1000 ;
	    RECT 109.1000 80.8000 109.5000 83.1000 ;
	    RECT 110.2000 80.8000 110.6000 83.1000 ;
	    RECT 111.8000 80.8000 112.2000 84.9000 ;
	    RECT 113.4000 80.8000 113.8000 85.1000 ;
	    RECT 116.6000 80.8000 117.0000 85.1000 ;
	    RECT 118.2000 80.8000 118.6000 82.9000 ;
	    RECT 119.8000 80.8000 120.2000 83.1000 ;
	    RECT 120.6000 80.8000 121.0000 85.1000 ;
	    RECT 122.2000 80.8000 122.6000 85.1000 ;
	    RECT 123.8000 80.8000 124.2000 85.1000 ;
	    RECT 126.6000 80.8000 127.0000 83.1000 ;
	    RECT 128.2000 80.8000 128.6000 83.1000 ;
	    RECT 131.0000 80.8000 131.4000 85.0000 ;
	    RECT 133.4000 80.8000 133.8000 85.0000 ;
	    RECT 136.2000 80.8000 136.6000 83.1000 ;
	    RECT 137.8000 80.8000 138.2000 83.1000 ;
	    RECT 140.6000 80.8000 141.0000 85.1000 ;
	    RECT 142.2000 80.8000 142.6000 85.1000 ;
	    RECT 143.8000 80.8000 144.2000 84.5000 ;
	    RECT 146.2000 80.8000 146.6000 84.5000 ;
	    RECT 0.2000 80.2000 148.6000 80.8000 ;
	    RECT 1.4000 76.5000 1.8000 80.2000 ;
	    RECT 7.8000 76.9000 8.2000 80.2000 ;
	    RECT 9.4000 77.9000 9.8000 80.2000 ;
	    RECT 11.0000 76.1000 11.4000 80.2000 ;
	    RECT 12.6000 77.9000 13.0000 80.2000 ;
	    RECT 14.2000 76.1000 14.6000 80.2000 ;
	    RECT 15.8000 77.9000 16.2000 80.2000 ;
	    RECT 17.4000 77.9000 17.8000 80.2000 ;
	    RECT 19.0000 78.1000 19.4000 80.2000 ;
	    RECT 20.6000 77.9000 21.0000 80.2000 ;
	    RECT 22.5000 75.9000 22.9000 80.2000 ;
	    RECT 24.6000 77.9000 25.0000 80.2000 ;
	    RECT 26.2000 77.9000 26.6000 80.2000 ;
	    RECT 27.0000 75.9000 27.4000 80.2000 ;
	    RECT 28.6000 76.5000 29.0000 80.2000 ;
	    RECT 30.2000 75.9000 30.6000 80.2000 ;
	    RECT 32.6000 75.9000 33.0000 80.2000 ;
	    RECT 36.1000 75.9000 36.5000 80.2000 ;
	    RECT 39.8000 75.9000 40.2000 80.2000 ;
	    RECT 40.6000 77.9000 41.0000 80.2000 ;
	    RECT 42.2000 77.9000 42.6000 80.2000 ;
	    RECT 44.6000 75.9000 45.0000 80.2000 ;
	    RECT 45.4000 77.9000 45.8000 80.2000 ;
	    RECT 47.0000 77.9000 47.4000 80.2000 ;
	    RECT 49.4000 77.9000 49.8000 80.2000 ;
	    RECT 51.8000 76.5000 52.2000 80.2000 ;
	    RECT 55.8000 76.5000 56.2000 80.2000 ;
	    RECT 57.4000 75.9000 57.8000 80.2000 ;
	    RECT 59.0000 75.9000 59.4000 80.2000 ;
	    RECT 60.6000 75.9000 61.0000 80.2000 ;
	    RECT 62.2000 75.9000 62.6000 80.2000 ;
	    RECT 65.0000 77.9000 65.4000 80.2000 ;
	    RECT 66.6000 77.9000 67.0000 80.2000 ;
	    RECT 69.4000 76.0000 69.8000 80.2000 ;
	    RECT 71.8000 76.6000 72.3000 80.2000 ;
	    RECT 74.9000 79.9000 75.3000 80.2000 ;
	    RECT 74.9000 76.6000 75.4000 79.9000 ;
	    RECT 78.2000 75.9000 78.6000 80.2000 ;
	    RECT 79.0000 77.9000 79.4000 80.2000 ;
	    RECT 80.6000 77.9000 81.0000 80.2000 ;
	    RECT 82.2000 76.1000 82.6000 80.2000 ;
	    RECT 83.8000 77.9000 84.2000 80.2000 ;
	    RECT 84.6000 77.9000 85.0000 80.2000 ;
	    RECT 86.2000 78.1000 86.6000 80.2000 ;
	    RECT 88.6000 78.1000 89.0000 80.2000 ;
	    RECT 90.2000 77.9000 90.6000 80.2000 ;
	    RECT 91.8000 76.1000 92.2000 80.2000 ;
	    RECT 94.4000 75.9000 94.8000 80.2000 ;
	    RECT 95.8000 77.9000 96.2000 80.2000 ;
	    RECT 97.4000 78.1000 97.8000 80.2000 ;
	    RECT 105.4000 76.9000 105.8000 80.2000 ;
	    RECT 107.8000 78.1000 108.2000 80.2000 ;
	    RECT 109.4000 77.9000 109.8000 80.2000 ;
	    RECT 110.2000 75.9000 110.6000 80.2000 ;
	    RECT 112.3000 77.9000 112.7000 80.2000 ;
	    RECT 113.4000 75.9000 113.8000 80.2000 ;
	    RECT 115.5000 77.9000 115.9000 80.2000 ;
	    RECT 118.2000 76.5000 118.6000 80.2000 ;
	    RECT 119.8000 77.9000 120.2000 80.2000 ;
	    RECT 121.4000 76.1000 121.8000 80.2000 ;
	    RECT 123.0000 75.9000 123.4000 80.2000 ;
	    RECT 125.1000 77.9000 125.5000 80.2000 ;
	    RECT 126.2000 77.9000 126.6000 80.2000 ;
	    RECT 127.8000 76.1000 128.2000 80.2000 ;
	    RECT 129.4000 75.9000 129.8000 80.2000 ;
	    RECT 131.5000 77.9000 131.9000 80.2000 ;
	    RECT 132.6000 75.9000 133.0000 80.2000 ;
	    RECT 134.2000 75.9000 134.6000 80.2000 ;
	    RECT 136.3000 77.9000 136.7000 80.2000 ;
	    RECT 137.4000 75.9000 137.8000 80.2000 ;
	    RECT 139.5000 77.9000 139.9000 80.2000 ;
	    RECT 142.2000 76.5000 142.6000 80.2000 ;
	    RECT 144.6000 76.5000 145.0000 80.2000 ;
	    RECT 1.4000 60.8000 1.8000 64.5000 ;
	    RECT 3.8000 60.8000 4.2000 65.1000 ;
	    RECT 6.6000 60.8000 7.0000 63.1000 ;
	    RECT 8.2000 60.8000 8.6000 63.1000 ;
	    RECT 11.0000 60.8000 11.4000 65.0000 ;
	    RECT 12.6000 60.8000 13.0000 65.1000 ;
	    RECT 15.0000 60.8000 15.5000 64.4000 ;
	    RECT 18.1000 61.1000 18.6000 64.4000 ;
	    RECT 18.1000 60.8000 18.5000 61.1000 ;
	    RECT 20.6000 60.8000 21.0000 64.5000 ;
	    RECT 23.3000 60.8000 23.7000 63.1000 ;
	    RECT 25.4000 60.8000 25.8000 65.1000 ;
	    RECT 27.0000 60.8000 27.4000 62.9000 ;
	    RECT 28.6000 60.8000 29.0000 63.1000 ;
	    RECT 29.7000 60.8000 30.1000 63.1000 ;
	    RECT 31.8000 60.8000 32.2000 65.1000 ;
	    RECT 32.6000 60.8000 33.0000 63.1000 ;
	    RECT 34.2000 60.8000 34.6000 62.9000 ;
	    RECT 36.1000 60.8000 36.5000 63.1000 ;
	    RECT 38.2000 60.8000 38.6000 65.1000 ;
	    RECT 39.8000 60.8000 40.2000 63.1000 ;
	    RECT 40.6000 60.8000 41.0000 63.1000 ;
	    RECT 42.2000 60.8000 42.6000 63.1000 ;
	    RECT 43.0000 60.8000 43.4000 63.1000 ;
	    RECT 44.6000 60.8000 45.0000 63.1000 ;
	    RECT 47.0000 60.8000 47.4000 64.5000 ;
	    RECT 55.0000 60.8000 55.4000 64.1000 ;
	    RECT 56.6000 60.8000 57.0000 65.1000 ;
	    RECT 58.7000 60.8000 59.1000 63.1000 ;
	    RECT 59.8000 60.8000 60.2000 63.1000 ;
	    RECT 61.4000 60.8000 61.8000 63.1000 ;
	    RECT 62.2000 60.8000 62.6000 65.1000 ;
	    RECT 63.8000 60.8000 64.2000 64.5000 ;
	    RECT 66.2000 61.1000 66.7000 64.4000 ;
	    RECT 66.3000 60.8000 66.7000 61.1000 ;
	    RECT 69.3000 60.8000 69.8000 64.4000 ;
	    RECT 71.8000 60.8000 72.2000 64.5000 ;
	    RECT 73.4000 60.8000 73.8000 65.1000 ;
	    RECT 79.0000 60.8000 79.4000 64.1000 ;
	    RECT 82.2000 60.8000 82.6000 65.1000 ;
	    RECT 83.8000 60.8000 84.2000 64.9000 ;
	    RECT 85.4000 60.8000 85.8000 63.1000 ;
	    RECT 86.2000 60.8000 86.6000 63.1000 ;
	    RECT 87.8000 60.8000 88.2000 63.1000 ;
	    RECT 88.6000 60.8000 89.0000 63.1000 ;
	    RECT 90.2000 60.8000 90.6000 63.1000 ;
	    RECT 91.0000 60.8000 91.4000 65.1000 ;
	    RECT 94.2000 60.8000 94.6000 64.1000 ;
	    RECT 102.2000 60.8000 102.6000 64.9000 ;
	    RECT 103.8000 60.8000 104.2000 63.1000 ;
	    RECT 104.6000 60.8000 105.0000 63.1000 ;
	    RECT 106.2000 60.8000 106.6000 63.1000 ;
	    RECT 107.8000 60.8000 108.2000 62.9000 ;
	    RECT 109.4000 60.8000 109.8000 63.1000 ;
	    RECT 110.2000 60.8000 110.6000 65.1000 ;
	    RECT 112.3000 60.8000 112.7000 63.1000 ;
	    RECT 114.2000 60.8000 114.6000 62.9000 ;
	    RECT 115.8000 60.8000 116.2000 63.1000 ;
	    RECT 116.6000 60.8000 117.0000 65.1000 ;
	    RECT 119.0000 60.8000 119.4000 63.1000 ;
	    RECT 120.6000 60.8000 121.0000 62.9000 ;
	    RECT 122.2000 60.8000 122.6000 65.1000 ;
	    RECT 124.3000 60.8000 124.7000 63.1000 ;
	    RECT 126.2000 60.8000 126.6000 65.1000 ;
	    RECT 127.0000 60.8000 127.4000 65.1000 ;
	    RECT 129.1000 60.8000 129.5000 63.1000 ;
	    RECT 131.8000 60.8000 132.2000 64.5000 ;
	    RECT 133.7000 60.8000 134.1000 63.1000 ;
	    RECT 135.8000 60.8000 136.2000 65.1000 ;
	    RECT 136.6000 60.8000 137.0000 65.1000 ;
	    RECT 138.7000 60.8000 139.1000 63.1000 ;
	    RECT 140.6000 60.8000 141.0000 63.1000 ;
	    RECT 141.4000 60.8000 141.8000 63.1000 ;
	    RECT 143.0000 60.8000 143.4000 63.1000 ;
	    RECT 144.6000 60.8000 145.0000 63.1000 ;
	    RECT 146.2000 60.8000 146.6000 64.5000 ;
	    RECT 0.2000 60.2000 148.6000 60.8000 ;
	    RECT 1.4000 56.5000 1.8000 60.2000 ;
	    RECT 3.8000 56.5000 4.2000 60.2000 ;
	    RECT 5.4000 57.9000 5.8000 60.2000 ;
	    RECT 7.8000 56.5000 8.2000 60.2000 ;
	    RECT 10.2000 55.9000 10.6000 60.2000 ;
	    RECT 13.0000 57.9000 13.4000 60.2000 ;
	    RECT 14.6000 57.9000 15.0000 60.2000 ;
	    RECT 17.4000 56.0000 17.8000 60.2000 ;
	    RECT 19.9000 59.9000 20.3000 60.2000 ;
	    RECT 19.8000 56.6000 20.3000 59.9000 ;
	    RECT 22.9000 56.6000 23.4000 60.2000 ;
	    RECT 25.4000 56.0000 25.8000 60.2000 ;
	    RECT 28.2000 57.9000 28.6000 60.2000 ;
	    RECT 29.8000 57.9000 30.2000 60.2000 ;
	    RECT 32.6000 55.9000 33.0000 60.2000 ;
	    RECT 35.0000 56.5000 35.4000 60.2000 ;
	    RECT 36.6000 55.9000 37.0000 60.2000 ;
	    RECT 38.2000 56.5000 38.6000 60.2000 ;
	    RECT 39.8000 57.9000 40.2000 60.2000 ;
	    RECT 41.4000 57.9000 41.8000 60.2000 ;
	    RECT 43.0000 56.6000 43.5000 60.2000 ;
	    RECT 46.1000 59.9000 46.5000 60.2000 ;
	    RECT 50.3000 59.9000 50.7000 60.2000 ;
	    RECT 46.1000 56.6000 46.6000 59.9000 ;
	    RECT 50.2000 56.6000 50.7000 59.9000 ;
	    RECT 53.3000 56.6000 53.8000 60.2000 ;
	    RECT 55.8000 56.5000 56.2000 60.2000 ;
	    RECT 57.4000 55.9000 57.8000 60.2000 ;
	    RECT 59.0000 56.1000 59.4000 60.2000 ;
	    RECT 60.6000 57.9000 61.0000 60.2000 ;
	    RECT 61.4000 55.9000 61.8000 60.2000 ;
	    RECT 64.6000 57.9000 65.0000 60.2000 ;
	    RECT 65.4000 57.9000 65.8000 60.2000 ;
	    RECT 67.0000 57.9000 67.4000 60.2000 ;
	    RECT 67.8000 55.9000 68.2000 60.2000 ;
	    RECT 69.4000 56.5000 69.8000 60.2000 ;
	    RECT 71.0000 57.9000 71.4000 60.2000 ;
	    RECT 72.6000 57.9000 73.0000 60.2000 ;
	    RECT 73.4000 55.9000 73.8000 60.2000 ;
	    RECT 77.4000 55.9000 77.8000 60.2000 ;
	    RECT 78.2000 55.9000 78.6000 60.2000 ;
	    RECT 79.8000 56.5000 80.2000 60.2000 ;
	    RECT 81.4000 55.9000 81.8000 60.2000 ;
	    RECT 83.5000 57.9000 83.9000 60.2000 ;
	    RECT 84.6000 57.9000 85.0000 60.2000 ;
	    RECT 86.2000 57.9000 86.6000 60.2000 ;
	    RECT 87.0000 57.9000 87.4000 60.2000 ;
	    RECT 90.2000 55.9000 90.6000 60.2000 ;
	    RECT 93.4000 56.5000 93.8000 60.2000 ;
	    RECT 97.4000 55.9000 97.8000 60.2000 ;
	    RECT 100.2000 57.9000 100.6000 60.2000 ;
	    RECT 101.8000 57.9000 102.2000 60.2000 ;
	    RECT 104.6000 56.0000 105.0000 60.2000 ;
	    RECT 107.8000 55.9000 108.2000 60.2000 ;
	    RECT 109.4000 56.5000 109.8000 60.2000 ;
	    RECT 111.0000 55.9000 111.4000 60.2000 ;
	    RECT 112.1000 57.9000 112.5000 60.2000 ;
	    RECT 114.2000 55.9000 114.6000 60.2000 ;
	    RECT 115.0000 57.9000 115.4000 60.2000 ;
	    RECT 116.6000 56.1000 117.0000 60.2000 ;
	    RECT 118.2000 55.9000 118.6000 60.2000 ;
	    RECT 120.3000 57.9000 120.7000 60.2000 ;
	    RECT 121.7000 57.9000 122.1000 60.2000 ;
	    RECT 123.8000 55.9000 124.2000 60.2000 ;
	    RECT 124.6000 55.9000 125.0000 60.2000 ;
	    RECT 126.7000 57.9000 127.1000 60.2000 ;
	    RECT 127.8000 57.9000 128.2000 60.2000 ;
	    RECT 129.4000 57.9000 129.8000 60.2000 ;
	    RECT 131.0000 56.5000 131.4000 60.2000 ;
	    RECT 135.0000 56.5000 135.4000 60.2000 ;
	    RECT 137.4000 57.9000 137.8000 60.2000 ;
	    RECT 139.0000 56.5000 139.4000 60.2000 ;
	    RECT 140.6000 57.9000 141.0000 60.2000 ;
	    RECT 142.2000 57.9000 142.6000 60.2000 ;
	    RECT 143.8000 56.5000 144.2000 60.2000 ;
	    RECT 145.4000 57.9000 145.8000 60.2000 ;
	    RECT 147.0000 57.9000 147.4000 60.2000 ;
	    RECT 1.4000 40.8000 1.8000 45.1000 ;
	    RECT 4.2000 40.8000 4.6000 43.1000 ;
	    RECT 5.8000 40.8000 6.2000 43.1000 ;
	    RECT 8.6000 40.8000 9.0000 45.0000 ;
	    RECT 10.2000 40.8000 10.6000 45.1000 ;
	    RECT 13.4000 40.8000 13.8000 44.5000 ;
	    RECT 15.8000 40.8000 16.2000 44.5000 ;
	    RECT 17.4000 40.8000 17.8000 45.1000 ;
	    RECT 19.0000 40.8000 19.4000 44.5000 ;
	    RECT 21.4000 40.8000 21.8000 44.5000 ;
	    RECT 23.0000 40.8000 23.4000 45.1000 ;
	    RECT 24.6000 40.8000 25.0000 45.1000 ;
	    RECT 25.4000 40.8000 25.8000 43.1000 ;
	    RECT 27.8000 40.8000 28.2000 42.9000 ;
	    RECT 29.4000 40.8000 29.8000 43.1000 ;
	    RECT 30.2000 40.8000 30.6000 43.1000 ;
	    RECT 31.8000 40.8000 32.2000 44.9000 ;
	    RECT 33.4000 40.8000 33.8000 43.1000 ;
	    RECT 35.0000 40.8000 35.4000 42.9000 ;
	    RECT 37.4000 40.8000 37.8000 45.1000 ;
	    RECT 40.2000 40.8000 40.6000 43.1000 ;
	    RECT 41.8000 40.8000 42.2000 43.1000 ;
	    RECT 44.6000 40.8000 45.0000 45.0000 ;
	    RECT 48.6000 40.8000 49.0000 45.0000 ;
	    RECT 51.4000 40.8000 51.8000 43.1000 ;
	    RECT 53.0000 40.8000 53.4000 43.1000 ;
	    RECT 55.8000 40.8000 56.2000 45.1000 ;
	    RECT 58.2000 40.8000 58.6000 44.5000 ;
	    RECT 60.6000 40.8000 61.0000 44.5000 ;
	    RECT 62.2000 40.8000 62.6000 43.1000 ;
	    RECT 63.8000 40.8000 64.2000 43.1000 ;
	    RECT 65.4000 40.8000 65.8000 43.1000 ;
	    RECT 67.5000 40.8000 67.9000 45.1000 ;
	    RECT 69.4000 40.8000 69.8000 43.1000 ;
	    RECT 71.0000 40.8000 71.4000 43.1000 ;
	    RECT 72.6000 40.8000 73.0000 43.1000 ;
	    RECT 73.4000 40.8000 73.8000 45.1000 ;
	    RECT 77.4000 40.8000 77.8000 45.1000 ;
	    RECT 78.2000 40.8000 78.6000 43.1000 ;
	    RECT 79.8000 40.8000 80.2000 43.1000 ;
	    RECT 81.4000 40.8000 81.8000 45.1000 ;
	    RECT 82.2000 40.8000 82.6000 45.1000 ;
	    RECT 84.6000 40.8000 85.0000 43.1000 ;
	    RECT 86.2000 40.8000 86.6000 43.1000 ;
	    RECT 87.3000 40.8000 87.7000 43.1000 ;
	    RECT 89.4000 40.8000 89.8000 45.1000 ;
	    RECT 91.0000 40.8000 91.4000 44.5000 ;
	    RECT 94.5000 40.8000 94.9000 43.1000 ;
	    RECT 96.6000 40.8000 97.0000 45.1000 ;
	    RECT 98.2000 40.8000 98.6000 43.1000 ;
	    RECT 102.2000 40.8000 102.6000 45.1000 ;
	    RECT 103.8000 40.8000 104.2000 45.1000 ;
	    RECT 106.6000 40.8000 107.0000 43.1000 ;
	    RECT 108.2000 40.8000 108.6000 43.1000 ;
	    RECT 111.0000 40.8000 111.4000 45.0000 ;
	    RECT 112.6000 40.8000 113.0000 45.1000 ;
	    RECT 115.0000 40.8000 115.4000 44.5000 ;
	    RECT 116.6000 40.8000 117.0000 45.1000 ;
	    RECT 118.2000 40.8000 118.6000 45.0000 ;
	    RECT 121.0000 40.8000 121.4000 43.1000 ;
	    RECT 122.6000 40.8000 123.0000 43.1000 ;
	    RECT 125.4000 40.8000 125.8000 45.1000 ;
	    RECT 127.8000 40.8000 128.2000 44.5000 ;
	    RECT 130.2000 40.8000 130.6000 45.1000 ;
	    RECT 132.9000 40.8000 133.3000 43.1000 ;
	    RECT 135.0000 40.8000 135.4000 45.1000 ;
	    RECT 135.8000 40.8000 136.2000 43.1000 ;
	    RECT 137.4000 40.8000 137.8000 45.1000 ;
	    RECT 139.5000 40.8000 139.9000 43.1000 ;
	    RECT 141.4000 40.8000 141.8000 44.5000 ;
	    RECT 143.8000 40.8000 144.2000 44.5000 ;
	    RECT 146.2000 40.8000 146.6000 43.1000 ;
	    RECT 0.2000 40.2000 148.6000 40.8000 ;
	    RECT 1.4000 36.5000 1.8000 40.2000 ;
	    RECT 3.8000 35.9000 4.2000 40.2000 ;
	    RECT 6.6000 37.9000 7.0000 40.2000 ;
	    RECT 8.2000 37.9000 8.6000 40.2000 ;
	    RECT 11.0000 36.0000 11.4000 40.2000 ;
	    RECT 12.6000 37.9000 13.0000 40.2000 ;
	    RECT 14.2000 35.9000 14.6000 40.2000 ;
	    RECT 16.6000 37.9000 17.0000 40.2000 ;
	    RECT 18.2000 37.9000 18.6000 40.2000 ;
	    RECT 19.0000 37.9000 19.4000 40.2000 ;
	    RECT 20.6000 37.9000 21.0000 40.2000 ;
	    RECT 22.2000 38.1000 22.6000 40.2000 ;
	    RECT 23.8000 37.9000 24.2000 40.2000 ;
	    RECT 29.4000 36.9000 29.8000 40.2000 ;
	    RECT 31.0000 35.9000 31.4000 40.2000 ;
	    RECT 35.0000 35.9000 35.4000 40.2000 ;
	    RECT 36.6000 37.9000 37.0000 40.2000 ;
	    RECT 37.4000 35.9000 37.8000 40.2000 ;
	    RECT 39.5000 37.9000 39.9000 40.2000 ;
	    RECT 41.7000 35.9000 42.1000 40.2000 ;
	    RECT 43.8000 37.9000 44.2000 40.2000 ;
	    RECT 45.4000 37.9000 45.8000 40.2000 ;
	    RECT 46.2000 37.9000 46.6000 40.2000 ;
	    RECT 49.7000 37.9000 50.1000 40.2000 ;
	    RECT 51.8000 35.9000 52.2000 40.2000 ;
	    RECT 52.9000 37.9000 53.3000 40.2000 ;
	    RECT 55.0000 35.9000 55.4000 40.2000 ;
	    RECT 55.8000 35.9000 56.2000 40.2000 ;
	    RECT 58.5000 37.9000 58.9000 40.2000 ;
	    RECT 60.6000 35.9000 61.0000 40.2000 ;
	    RECT 61.4000 35.9000 61.8000 40.2000 ;
	    RECT 63.0000 35.9000 63.4000 40.2000 ;
	    RECT 63.8000 37.9000 64.2000 40.2000 ;
	    RECT 65.4000 37.9000 65.8000 40.2000 ;
	    RECT 67.0000 36.9000 67.4000 40.2000 ;
	    RECT 72.6000 37.9000 73.0000 40.2000 ;
	    RECT 74.2000 37.9000 74.6000 40.2000 ;
	    RECT 75.0000 37.9000 75.4000 40.2000 ;
	    RECT 76.6000 38.1000 77.0000 40.2000 ;
	    RECT 78.2000 37.9000 78.6000 40.2000 ;
	    RECT 80.6000 36.5000 81.0000 40.2000 ;
	    RECT 83.0000 35.9000 83.4000 40.2000 ;
	    RECT 85.4000 37.9000 85.8000 40.2000 ;
	    RECT 87.0000 37.9000 87.4000 40.2000 ;
	    RECT 89.4000 35.9000 89.8000 40.2000 ;
	    RECT 91.8000 35.9000 92.2000 40.2000 ;
	    RECT 93.4000 37.9000 93.8000 40.2000 ;
	    RECT 94.2000 35.9000 94.6000 40.2000 ;
	    RECT 95.8000 36.5000 96.2000 40.2000 ;
	    RECT 99.0000 35.9000 99.4000 40.2000 ;
	    RECT 100.6000 36.5000 101.0000 40.2000 ;
	    RECT 102.2000 35.9000 102.6000 40.2000 ;
	    RECT 104.3000 37.9000 104.7000 40.2000 ;
	    RECT 105.4000 37.9000 105.8000 40.2000 ;
	    RECT 107.0000 36.1000 107.4000 40.2000 ;
	    RECT 108.6000 35.9000 109.0000 40.2000 ;
	    RECT 110.7000 37.9000 111.1000 40.2000 ;
	    RECT 112.6000 36.0000 113.0000 40.2000 ;
	    RECT 115.4000 37.9000 115.8000 40.2000 ;
	    RECT 117.0000 37.9000 117.4000 40.2000 ;
	    RECT 119.8000 35.9000 120.2000 40.2000 ;
	    RECT 122.2000 36.5000 122.6000 40.2000 ;
	    RECT 125.4000 36.0000 125.8000 40.2000 ;
	    RECT 128.2000 37.9000 128.6000 40.2000 ;
	    RECT 129.8000 37.9000 130.2000 40.2000 ;
	    RECT 132.6000 35.9000 133.0000 40.2000 ;
	    RECT 135.0000 36.5000 135.4000 40.2000 ;
	    RECT 139.0000 35.9000 139.4000 40.2000 ;
	    RECT 140.6000 37.9000 141.0000 40.2000 ;
	    RECT 142.2000 36.5000 142.6000 40.2000 ;
	    RECT 144.6000 36.5000 145.0000 40.2000 ;
	    RECT 1.4000 20.8000 1.8000 25.1000 ;
	    RECT 4.2000 20.8000 4.6000 23.1000 ;
	    RECT 5.8000 20.8000 6.2000 23.1000 ;
	    RECT 8.6000 20.8000 9.0000 25.0000 ;
	    RECT 10.5000 20.8000 10.9000 23.1000 ;
	    RECT 12.6000 20.8000 13.0000 25.1000 ;
	    RECT 13.4000 20.8000 13.8000 23.1000 ;
	    RECT 15.0000 20.8000 15.4000 23.1000 ;
	    RECT 20.6000 20.8000 21.0000 24.1000 ;
	    RECT 22.2000 20.8000 22.6000 25.1000 ;
	    RECT 24.3000 20.8000 24.7000 23.1000 ;
	    RECT 27.0000 20.8000 27.4000 25.1000 ;
	    RECT 32.6000 20.8000 33.0000 24.1000 ;
	    RECT 35.8000 20.8000 36.2000 25.1000 ;
	    RECT 37.4000 20.8000 37.8000 24.5000 ;
	    RECT 39.8000 20.8000 40.2000 25.1000 ;
	    RECT 43.0000 20.8000 43.4000 25.1000 ;
	    RECT 45.4000 20.8000 45.8000 25.1000 ;
	    RECT 47.8000 20.8000 48.2000 25.1000 ;
	    RECT 51.0000 20.8000 51.4000 25.1000 ;
	    RECT 53.4000 20.8000 53.8000 25.1000 ;
	    RECT 55.0000 20.8000 55.4000 22.9000 ;
	    RECT 56.6000 20.8000 57.0000 23.1000 ;
	    RECT 57.7000 20.8000 58.1000 23.1000 ;
	    RECT 59.8000 20.8000 60.2000 25.1000 ;
	    RECT 62.2000 20.8000 62.6000 25.1000 ;
	    RECT 63.8000 20.8000 64.2000 22.9000 ;
	    RECT 65.4000 20.8000 65.8000 23.1000 ;
	    RECT 67.0000 20.8000 67.4000 24.1000 ;
	    RECT 72.6000 20.8000 73.0000 25.1000 ;
	    RECT 74.5000 20.8000 74.9000 23.1000 ;
	    RECT 76.6000 20.8000 77.0000 25.1000 ;
	    RECT 79.0000 20.8000 79.4000 25.1000 ;
	    RECT 79.8000 20.8000 80.2000 23.1000 ;
	    RECT 81.4000 20.8000 81.8000 24.9000 ;
	    RECT 83.8000 20.8000 84.2000 23.1000 ;
	    RECT 84.6000 20.8000 85.0000 23.1000 ;
	    RECT 86.2000 20.8000 86.6000 23.1000 ;
	    RECT 87.0000 20.8000 87.4000 25.1000 ;
	    RECT 89.4000 20.8000 89.8000 25.0000 ;
	    RECT 92.2000 20.8000 92.6000 23.1000 ;
	    RECT 93.8000 20.8000 94.2000 23.1000 ;
	    RECT 96.6000 20.8000 97.0000 25.1000 ;
	    RECT 100.6000 20.8000 101.0000 24.5000 ;
	    RECT 103.0000 20.8000 103.4000 24.5000 ;
	    RECT 105.4000 20.8000 105.8000 25.1000 ;
	    RECT 108.2000 20.8000 108.6000 23.1000 ;
	    RECT 109.8000 20.8000 110.2000 23.1000 ;
	    RECT 112.6000 20.8000 113.0000 25.0000 ;
	    RECT 114.2000 20.8000 114.6000 23.1000 ;
	    RECT 115.8000 20.8000 116.2000 25.1000 ;
	    RECT 119.0000 20.8000 119.4000 25.0000 ;
	    RECT 121.8000 20.8000 122.2000 23.1000 ;
	    RECT 123.4000 20.8000 123.8000 23.1000 ;
	    RECT 126.2000 20.8000 126.6000 25.1000 ;
	    RECT 129.4000 20.8000 129.8000 25.1000 ;
	    RECT 131.0000 20.8000 131.4000 24.5000 ;
	    RECT 135.0000 20.8000 135.4000 25.1000 ;
	    RECT 136.6000 20.8000 137.0000 25.0000 ;
	    RECT 139.4000 20.8000 139.8000 23.1000 ;
	    RECT 141.0000 20.8000 141.4000 23.1000 ;
	    RECT 143.8000 20.8000 144.2000 25.1000 ;
	    RECT 146.2000 20.8000 146.6000 24.5000 ;
	    RECT 0.2000 20.2000 148.6000 20.8000 ;
	    RECT 1.4000 15.9000 1.8000 20.2000 ;
	    RECT 4.2000 17.9000 4.6000 20.2000 ;
	    RECT 5.8000 19.2000 6.2000 20.2000 ;
	    RECT 5.8000 18.8000 6.6000 19.2000 ;
	    RECT 5.8000 17.9000 6.2000 18.8000 ;
	    RECT 8.6000 16.0000 9.0000 20.2000 ;
	    RECT 11.0000 15.9000 11.4000 20.2000 ;
	    RECT 13.8000 17.9000 14.2000 20.2000 ;
	    RECT 15.4000 17.9000 15.8000 20.2000 ;
	    RECT 18.2000 16.0000 18.6000 20.2000 ;
	    RECT 20.6000 18.1000 21.0000 20.2000 ;
	    RECT 22.2000 17.9000 22.6000 20.2000 ;
	    RECT 23.8000 17.9000 24.2000 20.2000 ;
	    RECT 24.6000 17.9000 25.0000 20.2000 ;
	    RECT 26.2000 18.1000 26.6000 20.2000 ;
	    RECT 27.8000 15.9000 28.2000 20.2000 ;
	    RECT 30.2000 17.9000 30.6000 20.2000 ;
	    RECT 31.8000 17.9000 32.2000 20.2000 ;
	    RECT 32.9000 17.9000 33.3000 20.2000 ;
	    RECT 35.0000 15.9000 35.4000 20.2000 ;
	    RECT 35.8000 15.9000 36.2000 20.2000 ;
	    RECT 39.0000 17.9000 39.4000 20.2000 ;
	    RECT 39.8000 17.9000 40.2000 20.2000 ;
	    RECT 41.4000 17.9000 41.8000 20.2000 ;
	    RECT 42.2000 17.9000 42.6000 20.2000 ;
	    RECT 43.8000 18.1000 44.2000 20.2000 ;
	    RECT 47.0000 15.9000 47.4000 20.2000 ;
	    RECT 49.4000 15.9000 49.8000 20.2000 ;
	    RECT 52.6000 15.9000 53.0000 20.2000 ;
	    RECT 53.7000 17.9000 54.1000 20.2000 ;
	    RECT 55.8000 15.9000 56.2000 20.2000 ;
	    RECT 56.6000 15.9000 57.0000 20.2000 ;
	    RECT 59.0000 16.5000 59.4000 20.2000 ;
	    RECT 63.0000 15.9000 63.4000 20.2000 ;
	    RECT 63.8000 17.9000 64.2000 20.2000 ;
	    RECT 65.4000 17.9000 65.8000 20.2000 ;
	    RECT 67.8000 15.9000 68.2000 20.2000 ;
	    RECT 68.6000 17.9000 69.0000 20.2000 ;
	    RECT 70.2000 17.9000 70.6000 20.2000 ;
	    RECT 71.8000 17.9000 72.2000 20.2000 ;
	    RECT 73.4000 16.9000 73.8000 20.2000 ;
	    RECT 79.8000 16.9000 80.2000 20.2000 ;
	    RECT 86.2000 16.9000 86.6000 20.2000 ;
	    RECT 93.4000 15.9000 93.8000 20.2000 ;
	    RECT 95.8000 15.9000 96.2000 20.2000 ;
	    RECT 96.6000 17.9000 97.0000 20.2000 ;
	    RECT 98.2000 17.9000 98.6000 20.2000 ;
	    RECT 101.4000 16.5000 101.8000 20.2000 ;
	    RECT 103.8000 15.9000 104.2000 20.2000 ;
	    RECT 106.2000 15.9000 106.6000 20.2000 ;
	    RECT 110.2000 16.5000 110.6000 20.2000 ;
	    RECT 111.8000 15.9000 112.2000 20.2000 ;
	    RECT 113.4000 16.5000 113.8000 20.2000 ;
	    RECT 115.8000 16.5000 116.2000 20.2000 ;
	    RECT 117.4000 15.9000 117.8000 20.2000 ;
	    RECT 118.2000 15.9000 118.6000 20.2000 ;
	    RECT 119.8000 16.5000 120.2000 20.2000 ;
	    RECT 123.0000 15.9000 123.4000 20.2000 ;
	    RECT 124.6000 17.9000 125.0000 20.2000 ;
	    RECT 126.2000 15.9000 126.6000 20.2000 ;
	    RECT 129.0000 17.9000 129.4000 20.2000 ;
	    RECT 130.6000 17.9000 131.0000 20.2000 ;
	    RECT 133.4000 16.0000 133.8000 20.2000 ;
	    RECT 135.8000 16.0000 136.2000 20.2000 ;
	    RECT 138.6000 17.9000 139.0000 20.2000 ;
	    RECT 140.2000 17.9000 140.6000 20.2000 ;
	    RECT 143.0000 15.9000 143.4000 20.2000 ;
	    RECT 145.4000 16.5000 145.8000 20.2000 ;
	    RECT 147.0000 15.9000 147.4000 20.2000 ;
	    RECT 6.2000 15.1000 6.6000 15.2000 ;
	    RECT 6.2000 14.8000 8.7000 15.1000 ;
	    RECT 8.3000 14.7000 8.7000 14.8000 ;
	    RECT 1.4000 0.8000 1.8000 4.5000 ;
	    RECT 3.0000 0.8000 3.4000 5.1000 ;
	    RECT 5.4000 0.8000 5.8000 4.5000 ;
	    RECT 7.8000 0.8000 8.2000 5.1000 ;
	    RECT 10.2000 0.8000 10.6000 3.1000 ;
	    RECT 11.8000 0.8000 12.2000 3.1000 ;
	    RECT 17.4000 0.8000 17.8000 4.1000 ;
	    RECT 20.6000 0.8000 21.0000 5.1000 ;
	    RECT 22.2000 0.8000 22.6000 4.1000 ;
	    RECT 27.8000 0.8000 28.2000 5.1000 ;
	    RECT 29.4000 0.8000 29.8000 5.1000 ;
	    RECT 31.5000 0.8000 31.9000 3.1000 ;
	    RECT 32.9000 0.8000 33.3000 3.1000 ;
	    RECT 35.0000 0.8000 35.4000 5.1000 ;
	    RECT 36.6000 0.8000 37.0000 4.1000 ;
	    RECT 42.2000 0.8000 42.6000 3.1000 ;
	    RECT 43.8000 0.8000 44.2000 2.9000 ;
	    RECT 47.0000 0.8000 47.4000 5.1000 ;
	    RECT 49.4000 0.8000 49.8000 5.1000 ;
	    RECT 51.5000 0.8000 51.9000 3.1000 ;
	    RECT 53.4000 0.8000 53.8000 4.1000 ;
	    RECT 59.0000 0.8000 59.4000 5.1000 ;
	    RECT 61.1000 0.8000 61.5000 3.1000 ;
	    RECT 62.2000 0.8000 62.6000 3.1000 ;
	    RECT 63.8000 0.8000 64.2000 3.1000 ;
	    RECT 65.4000 0.8000 65.8000 4.5000 ;
	    RECT 67.0000 0.8000 67.4000 3.1000 ;
	    RECT 68.6000 0.8000 69.0000 2.9000 ;
	    RECT 71.0000 0.8000 71.4000 5.1000 ;
	    RECT 73.8000 0.8000 74.2000 3.1000 ;
	    RECT 75.4000 0.8000 75.8000 3.1000 ;
	    RECT 78.2000 0.8000 78.6000 5.0000 ;
	    RECT 80.6000 0.8000 81.0000 4.5000 ;
	    RECT 83.0000 0.8000 83.4000 4.5000 ;
	    RECT 85.4000 0.8000 85.8000 5.0000 ;
	    RECT 88.2000 0.8000 88.6000 3.1000 ;
	    RECT 89.8000 0.8000 90.2000 3.1000 ;
	    RECT 92.6000 0.8000 93.0000 5.1000 ;
	    RECT 95.0000 0.8000 95.4000 4.5000 ;
	    RECT 97.4000 0.8000 97.8000 4.5000 ;
	    RECT 101.4000 0.8000 101.8000 5.1000 ;
	    RECT 104.2000 0.8000 104.6000 3.1000 ;
	    RECT 105.8000 0.8000 106.2000 3.1000 ;
	    RECT 108.6000 0.8000 109.0000 5.0000 ;
	    RECT 111.0000 0.8000 111.4000 4.5000 ;
	    RECT 113.4000 0.8000 113.8000 4.5000 ;
	    RECT 115.8000 0.8000 116.2000 4.5000 ;
	    RECT 118.2000 0.8000 118.6000 4.5000 ;
	    RECT 120.6000 0.8000 121.0000 4.5000 ;
	    RECT 123.0000 0.8000 123.4000 4.5000 ;
	    RECT 125.4000 0.8000 125.8000 4.5000 ;
	    RECT 127.8000 1.1000 128.3000 4.4000 ;
	    RECT 127.9000 0.8000 128.3000 1.1000 ;
	    RECT 130.9000 0.8000 131.4000 4.4000 ;
	    RECT 133.4000 0.8000 133.8000 4.5000 ;
	    RECT 135.8000 0.8000 136.2000 4.5000 ;
	    RECT 138.2000 0.8000 138.6000 4.5000 ;
	    RECT 140.6000 0.8000 141.0000 4.5000 ;
	    RECT 143.0000 0.8000 143.4000 4.5000 ;
	    RECT 144.6000 0.8000 145.0000 3.1000 ;
	    RECT 146.2000 0.8000 146.6000 3.1000 ;
	    RECT 0.2000 0.2000 148.6000 0.8000 ;
         LAYER metal2 ;
	    RECT 47.2000 120.3000 48.8000 120.7000 ;
	    RECT 47.2000 100.3000 48.8000 100.7000 ;
	    RECT 47.2000 80.3000 48.8000 80.7000 ;
	    RECT 47.2000 60.3000 48.8000 60.7000 ;
	    RECT 47.2000 40.3000 48.8000 40.7000 ;
	    RECT 47.2000 20.3000 48.8000 20.7000 ;
	    RECT 6.2000 18.8000 6.6000 19.2000 ;
	    RECT 6.2000 15.2000 6.5000 18.8000 ;
	    RECT 6.2000 14.8000 6.6000 15.2000 ;
	    RECT 47.2000 0.3000 48.8000 0.7000 ;
         LAYER metal3 ;
	    RECT 47.2000 120.3000 48.8000 120.7000 ;
	    RECT 47.2000 100.3000 48.8000 100.7000 ;
	    RECT 47.2000 80.3000 48.8000 80.7000 ;
	    RECT 47.2000 60.3000 48.8000 60.7000 ;
	    RECT 47.2000 40.3000 48.8000 40.7000 ;
	    RECT 47.2000 20.3000 48.8000 20.7000 ;
	    RECT 47.2000 0.3000 48.8000 0.7000 ;
         LAYER metal4 ;
	    RECT 47.2000 120.3000 48.8000 120.7000 ;
	    RECT 47.2000 100.3000 48.8000 100.7000 ;
	    RECT 47.2000 80.3000 48.8000 80.7000 ;
	    RECT 47.2000 60.3000 48.8000 60.7000 ;
	    RECT 47.2000 40.3000 48.8000 40.7000 ;
	    RECT 47.2000 20.3000 48.8000 20.7000 ;
	    RECT 47.2000 0.3000 48.8000 0.7000 ;
         LAYER metal5 ;
	    RECT 47.2000 120.2000 48.8000 120.7000 ;
	    RECT 47.2000 100.2000 48.8000 100.7000 ;
	    RECT 47.2000 80.2000 48.8000 80.7000 ;
	    RECT 47.2000 60.2000 48.8000 60.7000 ;
	    RECT 47.2000 40.2000 48.8000 40.7000 ;
	    RECT 47.2000 20.2000 48.8000 20.7000 ;
	    RECT 47.2000 0.2000 48.8000 0.7000 ;
         LAYER metal6 ;
	    RECT 47.2000 -3.0000 48.8000 123.0000 ;
      END
   END vdd
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 1.4000 110.8000 1.8000 113.0000 ;
	    RECT 4.2000 110.8000 4.6000 112.1000 ;
	    RECT 5.8000 110.8000 6.3000 112.1000 ;
	    RECT 8.6000 110.8000 9.0000 113.1000 ;
	    RECT 11.0000 110.8000 11.4000 113.1000 ;
	    RECT 13.4000 110.8000 13.9000 112.8000 ;
	    RECT 16.5000 111.1000 17.0000 112.8000 ;
	    RECT 16.5000 110.8000 16.9000 111.1000 ;
	    RECT 18.2000 110.8000 18.6000 112.1000 ;
	    RECT 20.6000 110.8000 21.0000 113.1000 ;
	    RECT 23.0000 110.8000 23.4000 113.0000 ;
	    RECT 25.8000 110.8000 26.2000 112.1000 ;
	    RECT 27.4000 110.8000 27.9000 112.1000 ;
	    RECT 30.2000 110.8000 30.6000 113.1000 ;
	    RECT 32.6000 110.8000 33.1000 112.8000 ;
	    RECT 35.7000 111.1000 36.2000 112.8000 ;
	    RECT 35.7000 110.8000 36.1000 111.1000 ;
	    RECT 38.2000 110.8000 38.6000 112.7000 ;
	    RECT 40.9000 110.8000 41.3000 113.1000 ;
	    RECT 43.0000 110.8000 43.4000 112.1000 ;
	    RECT 43.8000 110.8000 44.2000 112.1000 ;
	    RECT 45.4000 110.8000 45.8000 112.1000 ;
	    RECT 47.0000 110.8000 47.4000 113.1000 ;
	    RECT 53.4000 110.8000 53.8000 111.9000 ;
	    RECT 55.0000 110.8000 55.4000 112.1000 ;
	    RECT 56.6000 110.8000 57.0000 112.1000 ;
	    RECT 58.2000 110.8000 58.6000 112.1000 ;
	    RECT 59.8000 111.1000 60.3000 112.8000 ;
	    RECT 59.9000 110.8000 60.3000 111.1000 ;
	    RECT 62.9000 110.8000 63.4000 112.8000 ;
	    RECT 66.2000 110.8000 66.6000 113.1000 ;
	    RECT 67.8000 110.8000 68.2000 113.1000 ;
	    RECT 69.4000 110.8000 69.8000 113.1000 ;
	    RECT 71.8000 110.8000 72.2000 113.1000 ;
	    RECT 74.5000 110.8000 75.0000 112.1000 ;
	    RECT 76.2000 110.8000 76.6000 112.1000 ;
	    RECT 79.0000 110.8000 79.4000 113.0000 ;
	    RECT 81.4000 110.8000 81.8000 113.1000 ;
	    RECT 83.8000 110.8000 84.2000 113.1000 ;
	    RECT 86.2000 110.8000 86.6000 113.1000 ;
	    RECT 88.6000 110.8000 89.0000 113.1000 ;
	    RECT 91.0000 110.8000 91.4000 113.1000 ;
	    RECT 93.4000 110.8000 93.8000 113.1000 ;
	    RECT 95.8000 111.1000 96.3000 112.8000 ;
	    RECT 95.9000 110.8000 96.3000 111.1000 ;
	    RECT 98.9000 110.8000 99.4000 112.8000 ;
	    RECT 103.0000 110.8000 103.4000 113.1000 ;
	    RECT 105.4000 110.8000 105.8000 113.1000 ;
	    RECT 107.0000 110.8000 107.4000 113.1000 ;
	    RECT 109.4000 110.8000 109.8000 113.1000 ;
	    RECT 112.6000 110.8000 113.0000 113.1000 ;
	    RECT 115.3000 110.8000 115.8000 112.1000 ;
	    RECT 117.0000 110.8000 117.4000 112.1000 ;
	    RECT 119.8000 110.8000 120.2000 113.0000 ;
	    RECT 122.2000 110.8000 122.6000 113.1000 ;
	    RECT 124.6000 110.8000 125.0000 113.1000 ;
	    RECT 127.0000 110.8000 127.4000 113.0000 ;
	    RECT 129.8000 110.8000 130.2000 112.1000 ;
	    RECT 131.4000 110.8000 131.9000 112.1000 ;
	    RECT 134.2000 110.8000 134.6000 113.1000 ;
	    RECT 136.6000 110.8000 137.0000 113.1000 ;
	    RECT 139.0000 110.8000 139.4000 113.1000 ;
	    RECT 141.4000 110.8000 141.8000 113.1000 ;
	    RECT 143.8000 110.8000 144.2000 113.1000 ;
	    RECT 146.2000 110.8000 146.6000 113.1000 ;
	    RECT 0.2000 110.2000 148.6000 110.8000 ;
	    RECT 1.4000 107.9000 1.8000 110.2000 ;
	    RECT 3.8000 108.0000 4.2000 110.2000 ;
	    RECT 6.6000 108.9000 7.0000 110.2000 ;
	    RECT 8.2000 108.9000 8.7000 110.2000 ;
	    RECT 11.0000 107.9000 11.4000 110.2000 ;
	    RECT 12.6000 108.9000 13.0000 110.2000 ;
	    RECT 14.2000 108.9000 14.6000 110.2000 ;
	    RECT 15.8000 108.9000 16.2000 110.2000 ;
	    RECT 17.4000 107.9000 17.8000 110.2000 ;
	    RECT 19.8000 108.0000 20.2000 110.2000 ;
	    RECT 22.6000 108.9000 23.0000 110.2000 ;
	    RECT 24.2000 108.9000 24.7000 110.2000 ;
	    RECT 27.0000 107.9000 27.4000 110.2000 ;
	    RECT 29.4000 108.2000 29.9000 110.2000 ;
	    RECT 32.5000 109.9000 32.9000 110.2000 ;
	    RECT 32.5000 108.2000 33.0000 109.9000 ;
	    RECT 37.4000 109.1000 37.8000 110.2000 ;
	    RECT 39.0000 108.9000 39.4000 110.2000 ;
	    RECT 40.6000 108.9000 41.0000 110.2000 ;
	    RECT 43.3000 108.0000 43.7000 110.2000 ;
	    RECT 47.0000 108.3000 47.4000 110.2000 ;
	    RECT 51.0000 108.9000 51.4000 110.2000 ;
	    RECT 52.6000 109.1000 53.0000 110.2000 ;
	    RECT 58.2000 108.3000 58.6000 110.2000 ;
	    RECT 61.4000 108.3000 61.8000 110.2000 ;
	    RECT 64.6000 107.9000 65.0000 110.2000 ;
	    RECT 65.4000 107.9000 65.8000 110.2000 ;
	    RECT 68.7000 109.9000 69.1000 110.2000 ;
	    RECT 68.6000 108.2000 69.1000 109.9000 ;
	    RECT 71.7000 108.2000 72.2000 110.2000 ;
	    RECT 74.2000 108.9000 74.6000 110.2000 ;
	    RECT 75.8000 108.0000 76.2000 110.2000 ;
	    RECT 78.6000 108.9000 79.0000 110.2000 ;
	    RECT 80.2000 108.9000 80.7000 110.2000 ;
	    RECT 83.0000 107.9000 83.4000 110.2000 ;
	    RECT 85.4000 107.9000 85.8000 110.2000 ;
	    RECT 87.8000 107.9000 88.2000 110.2000 ;
	    RECT 90.5000 108.9000 91.0000 110.2000 ;
	    RECT 92.2000 108.9000 92.6000 110.2000 ;
	    RECT 95.0000 108.0000 95.4000 110.2000 ;
	    RECT 99.0000 107.9000 99.4000 110.2000 ;
	    RECT 101.7000 108.9000 102.2000 110.2000 ;
	    RECT 103.4000 108.9000 103.8000 110.2000 ;
	    RECT 106.2000 108.0000 106.6000 110.2000 ;
	    RECT 107.8000 108.9000 108.2000 110.2000 ;
	    RECT 110.2000 107.7000 110.6000 110.2000 ;
	    RECT 112.8000 107.5000 113.2000 110.2000 ;
	    RECT 115.8000 108.3000 116.2000 110.2000 ;
	    RECT 118.2000 107.7000 118.6000 110.2000 ;
	    RECT 120.8000 107.5000 121.2000 110.2000 ;
	    RECT 122.5000 107.9000 122.9000 110.2000 ;
	    RECT 124.6000 108.9000 125.0000 110.2000 ;
	    RECT 125.4000 108.9000 125.8000 110.2000 ;
	    RECT 127.0000 108.9000 127.4000 110.2000 ;
	    RECT 128.6000 108.3000 129.0000 110.2000 ;
	    RECT 131.3000 107.9000 131.7000 110.2000 ;
	    RECT 133.4000 108.9000 133.8000 110.2000 ;
	    RECT 134.2000 108.9000 134.6000 110.2000 ;
	    RECT 135.8000 108.9000 136.2000 110.2000 ;
	    RECT 136.6000 108.9000 137.0000 110.2000 ;
	    RECT 138.2000 108.9000 138.6000 110.2000 ;
	    RECT 139.8000 107.9000 140.2000 110.2000 ;
	    RECT 142.5000 108.9000 143.0000 110.2000 ;
	    RECT 144.2000 108.9000 144.6000 110.2000 ;
	    RECT 147.0000 108.0000 147.4000 110.2000 ;
	    RECT 1.4000 90.8000 1.8000 93.1000 ;
	    RECT 3.8000 90.8000 4.2000 93.1000 ;
	    RECT 6.2000 90.8000 6.6000 93.0000 ;
	    RECT 9.0000 90.8000 9.4000 92.1000 ;
	    RECT 10.6000 90.8000 11.1000 92.1000 ;
	    RECT 13.4000 90.8000 13.8000 93.1000 ;
	    RECT 15.8000 90.8000 16.2000 93.0000 ;
	    RECT 18.6000 90.8000 19.0000 92.1000 ;
	    RECT 20.2000 90.8000 20.7000 92.1000 ;
	    RECT 23.0000 90.8000 23.4000 93.1000 ;
	    RECT 25.4000 90.8000 25.9000 92.8000 ;
	    RECT 28.5000 91.1000 29.0000 92.8000 ;
	    RECT 28.5000 90.8000 28.9000 91.1000 ;
	    RECT 31.0000 90.8000 31.4000 92.7000 ;
	    RECT 33.4000 90.8000 33.8000 92.1000 ;
	    RECT 35.0000 90.8000 35.4000 92.1000 ;
	    RECT 36.6000 90.8000 37.1000 92.8000 ;
	    RECT 39.7000 91.1000 40.2000 92.8000 ;
	    RECT 39.7000 90.8000 40.1000 91.1000 ;
	    RECT 41.4000 90.8000 41.8000 92.1000 ;
	    RECT 43.0000 90.8000 43.4000 92.1000 ;
	    RECT 44.6000 90.8000 45.0000 92.7000 ;
	    RECT 48.6000 90.8000 49.0000 92.1000 ;
	    RECT 50.7000 90.8000 51.1000 93.1000 ;
	    RECT 51.8000 90.8000 52.2000 92.1000 ;
	    RECT 53.9000 90.8000 54.3000 93.1000 ;
	    RECT 55.8000 90.8000 56.2000 92.1000 ;
	    RECT 56.6000 90.8000 57.0000 94.1000 ;
	    RECT 60.6000 90.8000 61.0000 93.1000 ;
	    RECT 62.5000 90.8000 62.9000 93.1000 ;
	    RECT 64.6000 90.8000 65.0000 92.1000 ;
	    RECT 67.0000 90.8000 67.4000 92.7000 ;
	    RECT 68.6000 90.8000 69.0000 92.1000 ;
	    RECT 70.2000 90.8000 70.6000 92.1000 ;
	    RECT 71.8000 90.8000 72.2000 92.1000 ;
	    RECT 73.4000 90.8000 73.8000 93.1000 ;
	    RECT 76.1000 90.8000 76.6000 92.1000 ;
	    RECT 77.8000 90.8000 78.2000 92.1000 ;
	    RECT 80.6000 90.8000 81.0000 93.0000 ;
	    RECT 83.0000 90.8000 83.4000 93.1000 ;
	    RECT 85.4000 90.8000 85.8000 93.1000 ;
	    RECT 87.6000 90.8000 88.0000 93.5000 ;
	    RECT 90.2000 90.8000 90.6000 93.3000 ;
	    RECT 92.6000 90.8000 93.0000 93.1000 ;
	    RECT 94.2000 90.8000 94.6000 92.1000 ;
	    RECT 95.8000 90.8000 96.2000 92.1000 ;
	    RECT 97.4000 90.8000 97.8000 93.1000 ;
	    RECT 100.6000 90.8000 101.0000 93.1000 ;
	    RECT 103.0000 90.8000 103.4000 93.0000 ;
	    RECT 105.8000 90.8000 106.2000 92.1000 ;
	    RECT 107.4000 90.8000 107.9000 92.1000 ;
	    RECT 110.2000 90.8000 110.6000 93.1000 ;
	    RECT 113.4000 90.8000 113.8000 92.7000 ;
	    RECT 116.6000 90.8000 117.0000 92.7000 ;
	    RECT 119.5000 90.8000 119.9000 93.0000 ;
	    RECT 122.2000 90.8000 122.6000 92.7000 ;
	    RECT 125.4000 90.8000 125.8000 92.7000 ;
	    RECT 128.6000 90.8000 129.0000 93.1000 ;
	    RECT 131.3000 90.8000 131.8000 92.1000 ;
	    RECT 133.0000 90.8000 133.4000 92.1000 ;
	    RECT 135.8000 90.8000 136.2000 93.0000 ;
	    RECT 137.4000 90.8000 137.8000 92.1000 ;
	    RECT 139.5000 90.8000 139.9000 93.1000 ;
	    RECT 141.4000 90.8000 141.8000 93.1000 ;
	    RECT 143.8000 90.8000 144.2000 92.1000 ;
	    RECT 145.4000 90.8000 145.8000 93.1000 ;
	    RECT 0.2000 90.2000 148.6000 90.8000 ;
	    RECT 1.4000 87.9000 1.8000 90.2000 ;
	    RECT 3.8000 88.0000 4.2000 90.2000 ;
	    RECT 6.6000 88.9000 7.0000 90.2000 ;
	    RECT 8.2000 88.9000 8.7000 90.2000 ;
	    RECT 11.0000 87.9000 11.4000 90.2000 ;
	    RECT 13.4000 88.2000 13.9000 90.2000 ;
	    RECT 16.5000 89.9000 16.9000 90.2000 ;
	    RECT 16.5000 88.2000 17.0000 89.9000 ;
	    RECT 19.0000 88.3000 19.4000 90.2000 ;
	    RECT 22.2000 87.9000 22.6000 90.2000 ;
	    RECT 23.8000 87.9000 24.2000 90.2000 ;
	    RECT 24.6000 88.9000 25.0000 90.2000 ;
	    RECT 26.2000 88.9000 26.6000 90.2000 ;
	    RECT 27.8000 88.9000 28.2000 90.2000 ;
	    RECT 29.4000 88.2000 29.9000 90.2000 ;
	    RECT 32.5000 89.9000 32.9000 90.2000 ;
	    RECT 32.5000 88.2000 33.0000 89.9000 ;
	    RECT 35.0000 87.9000 35.4000 90.2000 ;
	    RECT 37.7000 88.9000 38.2000 90.2000 ;
	    RECT 39.4000 88.9000 39.8000 90.2000 ;
	    RECT 42.2000 88.0000 42.6000 90.2000 ;
	    RECT 46.2000 86.9000 46.6000 90.2000 ;
	    RECT 50.2000 88.3000 50.6000 90.2000 ;
	    RECT 53.4000 88.3000 53.8000 90.2000 ;
	    RECT 55.8000 87.9000 56.2000 90.2000 ;
	    RECT 56.6000 88.9000 57.0000 90.2000 ;
	    RECT 60.6000 86.9000 61.0000 90.2000 ;
	    RECT 62.5000 88.0000 62.9000 90.2000 ;
	    RECT 65.4000 88.9000 65.8000 90.2000 ;
	    RECT 67.0000 88.3000 67.4000 90.2000 ;
	    RECT 69.4000 87.9000 69.8000 90.2000 ;
	    RECT 71.0000 87.9000 71.4000 90.2000 ;
	    RECT 73.5000 89.9000 73.9000 90.2000 ;
	    RECT 73.4000 88.2000 73.9000 89.9000 ;
	    RECT 76.5000 88.2000 77.0000 90.2000 ;
	    RECT 79.0000 88.0000 79.4000 90.2000 ;
	    RECT 81.8000 88.9000 82.2000 90.2000 ;
	    RECT 83.4000 88.9000 83.9000 90.2000 ;
	    RECT 86.2000 87.9000 86.6000 90.2000 ;
	    RECT 88.6000 87.9000 89.0000 90.2000 ;
	    RECT 90.2000 87.9000 90.6000 90.2000 ;
	    RECT 91.8000 87.9000 92.2000 90.2000 ;
	    RECT 94.2000 87.9000 94.6000 90.2000 ;
	    RECT 95.8000 87.9000 96.2000 90.2000 ;
	    RECT 98.2000 88.3000 98.6000 90.2000 ;
	    RECT 102.2000 87.9000 102.6000 90.2000 ;
	    RECT 103.8000 87.9000 104.2000 90.2000 ;
	    RECT 104.6000 87.9000 105.0000 90.2000 ;
	    RECT 106.2000 87.9000 106.6000 90.2000 ;
	    RECT 107.8000 88.3000 108.2000 90.2000 ;
	    RECT 111.5000 88.0000 111.9000 90.2000 ;
	    RECT 115.8000 88.3000 116.2000 90.2000 ;
	    RECT 119.8000 86.9000 120.2000 90.2000 ;
	    RECT 120.6000 87.9000 121.0000 90.2000 ;
	    RECT 122.2000 87.9000 122.6000 90.2000 ;
	    RECT 123.8000 88.0000 124.2000 90.2000 ;
	    RECT 126.6000 88.9000 127.0000 90.2000 ;
	    RECT 128.2000 88.9000 128.7000 90.2000 ;
	    RECT 131.0000 87.9000 131.4000 90.2000 ;
	    RECT 133.4000 87.9000 133.8000 90.2000 ;
	    RECT 136.1000 88.9000 136.6000 90.2000 ;
	    RECT 137.8000 88.9000 138.2000 90.2000 ;
	    RECT 140.6000 88.0000 141.0000 90.2000 ;
	    RECT 142.2000 87.9000 142.6000 90.2000 ;
	    RECT 143.8000 87.9000 144.2000 90.2000 ;
	    RECT 146.2000 87.9000 146.6000 90.2000 ;
	    RECT 1.4000 70.8000 1.8000 73.1000 ;
	    RECT 6.2000 70.8000 6.6000 71.9000 ;
	    RECT 7.8000 70.8000 8.2000 72.1000 ;
	    RECT 10.7000 70.8000 11.1000 73.0000 ;
	    RECT 13.9000 70.8000 14.3000 73.0000 ;
	    RECT 15.8000 70.8000 16.2000 73.1000 ;
	    RECT 20.6000 70.8000 21.0000 74.1000 ;
	    RECT 22.2000 70.8000 22.6000 72.9000 ;
	    RECT 23.8000 70.8000 24.2000 72.1000 ;
	    RECT 24.6000 70.8000 25.0000 73.1000 ;
	    RECT 27.0000 70.8000 27.4000 73.1000 ;
	    RECT 28.6000 70.8000 29.0000 73.1000 ;
	    RECT 30.2000 70.8000 30.6000 72.1000 ;
	    RECT 31.8000 70.8000 32.2000 72.1000 ;
	    RECT 32.6000 70.8000 33.0000 72.1000 ;
	    RECT 34.2000 70.8000 34.6000 72.1000 ;
	    RECT 35.8000 70.8000 36.2000 72.9000 ;
	    RECT 37.4000 70.8000 37.8000 72.1000 ;
	    RECT 38.2000 70.8000 38.6000 72.1000 ;
	    RECT 39.8000 70.8000 40.2000 72.1000 ;
	    RECT 42.2000 70.8000 42.6000 73.1000 ;
	    RECT 43.0000 70.8000 43.4000 72.1000 ;
	    RECT 44.6000 70.8000 45.0000 72.1000 ;
	    RECT 45.4000 70.8000 45.8000 73.1000 ;
	    RECT 49.4000 70.8000 49.8000 72.1000 ;
	    RECT 51.3000 70.8000 51.7000 73.1000 ;
	    RECT 53.4000 70.8000 53.8000 72.1000 ;
	    RECT 54.2000 70.8000 54.6000 72.1000 ;
	    RECT 56.3000 70.8000 56.7000 73.1000 ;
	    RECT 57.4000 70.8000 57.8000 73.1000 ;
	    RECT 59.0000 70.8000 59.4000 73.1000 ;
	    RECT 60.6000 70.8000 61.0000 73.1000 ;
	    RECT 62.2000 70.8000 62.6000 73.0000 ;
	    RECT 65.0000 70.8000 65.4000 72.1000 ;
	    RECT 66.6000 70.8000 67.1000 72.1000 ;
	    RECT 69.4000 70.8000 69.8000 73.1000 ;
	    RECT 71.8000 70.8000 72.3000 72.8000 ;
	    RECT 74.9000 71.1000 75.4000 72.8000 ;
	    RECT 74.9000 70.8000 75.3000 71.1000 ;
	    RECT 76.6000 70.8000 77.0000 72.1000 ;
	    RECT 78.2000 70.8000 78.6000 72.1000 ;
	    RECT 79.0000 70.8000 79.4000 73.1000 ;
	    RECT 82.5000 70.8000 82.9000 73.0000 ;
	    RECT 84.6000 70.8000 85.0000 74.1000 ;
	    RECT 90.2000 70.8000 90.6000 74.1000 ;
	    RECT 91.8000 70.8000 92.2000 73.3000 ;
	    RECT 94.4000 70.8000 94.8000 73.5000 ;
	    RECT 95.8000 70.8000 96.2000 74.1000 ;
	    RECT 103.8000 70.8000 104.2000 71.9000 ;
	    RECT 105.4000 70.8000 105.8000 72.1000 ;
	    RECT 109.4000 70.8000 109.8000 74.1000 ;
	    RECT 111.0000 70.8000 111.4000 72.7000 ;
	    RECT 114.2000 70.8000 114.6000 72.7000 ;
	    RECT 116.6000 70.8000 117.0000 72.1000 ;
	    RECT 118.7000 70.8000 119.1000 73.1000 ;
	    RECT 121.1000 70.8000 121.5000 73.0000 ;
	    RECT 123.8000 70.8000 124.2000 72.7000 ;
	    RECT 127.5000 70.8000 127.9000 73.0000 ;
	    RECT 130.2000 70.8000 130.6000 72.7000 ;
	    RECT 132.6000 70.8000 133.0000 73.1000 ;
	    RECT 135.0000 70.8000 135.4000 72.7000 ;
	    RECT 138.2000 70.8000 138.6000 72.7000 ;
	    RECT 140.6000 70.8000 141.0000 72.1000 ;
	    RECT 142.7000 70.8000 143.1000 73.1000 ;
	    RECT 144.6000 70.8000 145.0000 73.1000 ;
	    RECT 0.2000 70.2000 148.6000 70.8000 ;
	    RECT 1.4000 67.9000 1.8000 70.2000 ;
	    RECT 3.8000 68.0000 4.2000 70.2000 ;
	    RECT 6.6000 68.9000 7.0000 70.2000 ;
	    RECT 8.2000 68.9000 8.7000 70.2000 ;
	    RECT 11.0000 67.9000 11.4000 70.2000 ;
	    RECT 12.6000 67.9000 13.0000 70.2000 ;
	    RECT 15.0000 68.2000 15.5000 70.2000 ;
	    RECT 18.1000 69.9000 18.5000 70.2000 ;
	    RECT 18.1000 68.2000 18.6000 69.9000 ;
	    RECT 20.1000 67.9000 20.5000 70.2000 ;
	    RECT 22.2000 68.9000 22.6000 70.2000 ;
	    RECT 24.6000 68.3000 25.0000 70.2000 ;
	    RECT 28.6000 66.9000 29.0000 70.2000 ;
	    RECT 31.0000 68.3000 31.4000 70.2000 ;
	    RECT 32.6000 66.9000 33.0000 70.2000 ;
	    RECT 37.4000 68.3000 37.8000 70.2000 ;
	    RECT 39.8000 68.9000 40.2000 70.2000 ;
	    RECT 42.2000 67.9000 42.6000 70.2000 ;
	    RECT 43.0000 67.9000 43.4000 70.2000 ;
	    RECT 45.4000 68.9000 45.8000 70.2000 ;
	    RECT 47.5000 67.9000 47.9000 70.2000 ;
	    RECT 53.4000 69.1000 53.8000 70.2000 ;
	    RECT 55.0000 68.9000 55.4000 70.2000 ;
	    RECT 57.4000 68.3000 57.8000 70.2000 ;
	    RECT 59.8000 67.9000 60.2000 70.2000 ;
	    RECT 62.2000 67.9000 62.6000 70.2000 ;
	    RECT 63.8000 67.9000 64.2000 70.2000 ;
	    RECT 66.3000 69.9000 66.7000 70.2000 ;
	    RECT 66.2000 68.2000 66.7000 69.9000 ;
	    RECT 69.3000 68.2000 69.8000 70.2000 ;
	    RECT 71.8000 67.9000 72.2000 70.2000 ;
	    RECT 73.4000 67.9000 73.8000 70.2000 ;
	    RECT 77.4000 69.1000 77.8000 70.2000 ;
	    RECT 79.0000 68.9000 79.4000 70.2000 ;
	    RECT 80.6000 68.9000 81.0000 70.2000 ;
	    RECT 82.2000 68.9000 82.6000 70.2000 ;
	    RECT 84.1000 68.0000 84.5000 70.2000 ;
	    RECT 86.2000 67.9000 86.6000 70.2000 ;
	    RECT 88.6000 67.9000 89.0000 70.2000 ;
	    RECT 91.0000 68.9000 91.4000 70.2000 ;
	    RECT 92.6000 68.9000 93.0000 70.2000 ;
	    RECT 94.2000 68.9000 94.6000 70.2000 ;
	    RECT 95.8000 69.1000 96.2000 70.2000 ;
	    RECT 102.5000 68.0000 102.9000 70.2000 ;
	    RECT 106.2000 67.9000 106.6000 70.2000 ;
	    RECT 109.4000 66.9000 109.8000 70.2000 ;
	    RECT 111.0000 68.3000 111.4000 70.2000 ;
	    RECT 115.8000 66.9000 116.2000 70.2000 ;
	    RECT 116.6000 68.9000 117.0000 70.2000 ;
	    RECT 118.2000 68.9000 118.6000 70.2000 ;
	    RECT 119.0000 66.9000 119.4000 70.2000 ;
	    RECT 123.0000 68.3000 123.4000 70.2000 ;
	    RECT 126.2000 67.9000 126.6000 70.2000 ;
	    RECT 127.8000 68.3000 128.2000 70.2000 ;
	    RECT 130.2000 68.9000 130.6000 70.2000 ;
	    RECT 132.3000 67.9000 132.7000 70.2000 ;
	    RECT 135.0000 68.3000 135.4000 70.2000 ;
	    RECT 137.4000 68.3000 137.8000 70.2000 ;
	    RECT 140.6000 68.9000 141.0000 70.2000 ;
	    RECT 141.4000 67.9000 141.8000 70.2000 ;
	    RECT 144.6000 68.9000 145.0000 70.2000 ;
	    RECT 146.2000 67.9000 146.6000 70.2000 ;
	    RECT 1.4000 50.8000 1.8000 53.1000 ;
	    RECT 3.8000 50.8000 4.2000 53.1000 ;
	    RECT 5.4000 50.8000 5.8000 52.1000 ;
	    RECT 7.8000 50.8000 8.2000 53.1000 ;
	    RECT 10.2000 50.8000 10.6000 53.0000 ;
	    RECT 13.0000 50.8000 13.4000 52.1000 ;
	    RECT 14.6000 50.8000 15.1000 52.1000 ;
	    RECT 17.4000 50.8000 17.8000 53.1000 ;
	    RECT 19.8000 51.1000 20.3000 52.8000 ;
	    RECT 19.9000 50.8000 20.3000 51.1000 ;
	    RECT 22.9000 50.8000 23.4000 52.8000 ;
	    RECT 25.4000 50.8000 25.8000 53.1000 ;
	    RECT 28.1000 50.8000 28.6000 52.1000 ;
	    RECT 29.8000 50.8000 30.2000 52.1000 ;
	    RECT 32.6000 50.8000 33.0000 53.0000 ;
	    RECT 35.0000 50.8000 35.4000 53.1000 ;
	    RECT 36.6000 50.8000 37.0000 53.1000 ;
	    RECT 38.2000 50.8000 38.6000 53.1000 ;
	    RECT 41.4000 50.8000 41.8000 53.1000 ;
	    RECT 43.0000 50.8000 43.5000 52.8000 ;
	    RECT 46.1000 51.1000 46.6000 52.8000 ;
	    RECT 50.2000 51.1000 50.7000 52.8000 ;
	    RECT 46.1000 50.8000 46.5000 51.1000 ;
	    RECT 50.3000 50.8000 50.7000 51.1000 ;
	    RECT 53.3000 50.8000 53.8000 52.8000 ;
	    RECT 55.8000 50.8000 56.2000 53.1000 ;
	    RECT 57.4000 50.8000 57.8000 53.1000 ;
	    RECT 59.3000 50.8000 59.7000 53.0000 ;
	    RECT 61.4000 50.8000 61.8000 52.1000 ;
	    RECT 63.0000 50.8000 63.4000 52.1000 ;
	    RECT 64.6000 50.8000 65.0000 52.1000 ;
	    RECT 67.0000 50.8000 67.4000 53.1000 ;
	    RECT 67.8000 50.8000 68.2000 53.1000 ;
	    RECT 69.4000 50.8000 69.8000 53.1000 ;
	    RECT 71.0000 50.8000 71.4000 53.1000 ;
	    RECT 73.4000 50.8000 73.8000 52.1000 ;
	    RECT 75.0000 50.8000 75.4000 52.1000 ;
	    RECT 75.8000 50.8000 76.2000 52.1000 ;
	    RECT 77.4000 50.8000 77.8000 52.1000 ;
	    RECT 78.2000 50.8000 78.6000 53.1000 ;
	    RECT 79.8000 50.8000 80.2000 53.1000 ;
	    RECT 82.2000 50.8000 82.6000 52.7000 ;
	    RECT 86.2000 50.8000 86.6000 53.1000 ;
	    RECT 87.0000 50.8000 87.4000 52.1000 ;
	    RECT 88.6000 50.8000 89.0000 52.1000 ;
	    RECT 90.2000 50.8000 90.6000 52.1000 ;
	    RECT 91.0000 50.8000 91.4000 53.1000 ;
	    RECT 94.0000 50.8000 94.4000 53.1000 ;
	    RECT 97.4000 50.8000 97.8000 53.0000 ;
	    RECT 100.2000 50.8000 100.6000 52.1000 ;
	    RECT 101.8000 50.8000 102.3000 52.1000 ;
	    RECT 104.6000 50.8000 105.0000 53.1000 ;
	    RECT 106.2000 50.8000 106.6000 52.1000 ;
	    RECT 107.8000 50.8000 108.2000 52.1000 ;
	    RECT 109.4000 50.8000 109.8000 53.1000 ;
	    RECT 111.0000 50.8000 111.4000 53.1000 ;
	    RECT 113.4000 50.8000 113.8000 52.7000 ;
	    RECT 116.3000 50.8000 116.7000 53.0000 ;
	    RECT 119.0000 50.8000 119.4000 52.7000 ;
	    RECT 123.0000 50.8000 123.4000 52.7000 ;
	    RECT 125.4000 50.8000 125.8000 52.7000 ;
	    RECT 127.8000 50.8000 128.2000 53.1000 ;
	    RECT 130.5000 50.8000 130.9000 53.1000 ;
	    RECT 132.6000 50.8000 133.0000 52.1000 ;
	    RECT 133.4000 50.8000 133.8000 52.1000 ;
	    RECT 135.5000 50.8000 135.9000 53.1000 ;
	    RECT 137.4000 50.8000 137.8000 52.1000 ;
	    RECT 139.0000 50.8000 139.4000 53.1000 ;
	    RECT 140.6000 50.8000 141.0000 53.1000 ;
	    RECT 143.8000 50.8000 144.2000 53.1000 ;
	    RECT 145.4000 50.8000 145.8000 53.1000 ;
	    RECT 0.2000 50.2000 148.6000 50.8000 ;
	    RECT 1.4000 48.0000 1.8000 50.2000 ;
	    RECT 4.2000 48.9000 4.6000 50.2000 ;
	    RECT 5.8000 48.9000 6.3000 50.2000 ;
	    RECT 8.6000 47.9000 9.0000 50.2000 ;
	    RECT 10.2000 48.9000 10.6000 50.2000 ;
	    RECT 11.8000 48.9000 12.2000 50.2000 ;
	    RECT 13.4000 47.9000 13.8000 50.2000 ;
	    RECT 15.8000 47.9000 16.2000 50.2000 ;
	    RECT 17.4000 47.9000 17.8000 50.2000 ;
	    RECT 19.0000 47.9000 19.4000 50.2000 ;
	    RECT 21.4000 47.9000 21.8000 50.2000 ;
	    RECT 23.0000 47.9000 23.4000 50.2000 ;
	    RECT 24.6000 47.9000 25.0000 50.2000 ;
	    RECT 25.4000 48.9000 25.8000 50.2000 ;
	    RECT 29.4000 46.9000 29.8000 50.2000 ;
	    RECT 31.5000 48.0000 31.9000 50.2000 ;
	    RECT 33.4000 46.9000 33.8000 50.2000 ;
	    RECT 37.4000 48.0000 37.8000 50.2000 ;
	    RECT 40.2000 48.9000 40.6000 50.2000 ;
	    RECT 41.8000 48.9000 42.3000 50.2000 ;
	    RECT 44.6000 47.9000 45.0000 50.2000 ;
	    RECT 48.6000 47.9000 49.0000 50.2000 ;
	    RECT 51.3000 48.9000 51.8000 50.2000 ;
	    RECT 53.0000 48.9000 53.4000 50.2000 ;
	    RECT 55.8000 48.0000 56.2000 50.2000 ;
	    RECT 58.2000 47.9000 58.6000 50.2000 ;
	    RECT 60.6000 47.9000 61.0000 50.2000 ;
	    RECT 62.2000 48.9000 62.6000 50.2000 ;
	    RECT 65.4000 47.9000 65.8000 50.2000 ;
	    RECT 66.2000 48.9000 66.6000 50.2000 ;
	    RECT 67.8000 48.1000 68.2000 50.2000 ;
	    RECT 69.4000 47.9000 69.8000 50.2000 ;
	    RECT 72.6000 48.9000 73.0000 50.2000 ;
	    RECT 73.4000 48.9000 73.8000 50.2000 ;
	    RECT 75.0000 48.9000 75.4000 50.2000 ;
	    RECT 75.8000 48.9000 76.2000 50.2000 ;
	    RECT 77.4000 48.9000 77.8000 50.2000 ;
	    RECT 78.2000 47.9000 78.6000 50.2000 ;
	    RECT 81.4000 47.9000 81.8000 50.2000 ;
	    RECT 82.2000 48.9000 82.6000 50.2000 ;
	    RECT 83.8000 48.9000 84.2000 50.2000 ;
	    RECT 86.2000 47.9000 86.6000 50.2000 ;
	    RECT 88.6000 48.3000 89.0000 50.2000 ;
	    RECT 90.4000 47.9000 90.8000 50.2000 ;
	    RECT 93.4000 47.9000 93.8000 50.2000 ;
	    RECT 95.8000 48.3000 96.2000 50.2000 ;
	    RECT 98.2000 48.9000 98.6000 50.2000 ;
	    RECT 100.6000 48.9000 101.0000 50.2000 ;
	    RECT 102.2000 48.9000 102.6000 50.2000 ;
	    RECT 103.8000 48.0000 104.2000 50.2000 ;
	    RECT 106.6000 48.9000 107.0000 50.2000 ;
	    RECT 108.2000 48.9000 108.7000 50.2000 ;
	    RECT 111.0000 47.9000 111.4000 50.2000 ;
	    RECT 112.6000 47.9000 113.0000 50.2000 ;
	    RECT 115.0000 47.9000 115.4000 50.2000 ;
	    RECT 116.6000 47.9000 117.0000 50.2000 ;
	    RECT 118.2000 47.9000 118.6000 50.2000 ;
	    RECT 120.9000 48.9000 121.4000 50.2000 ;
	    RECT 122.6000 48.9000 123.0000 50.2000 ;
	    RECT 125.4000 48.0000 125.8000 50.2000 ;
	    RECT 127.3000 47.9000 127.7000 50.2000 ;
	    RECT 129.4000 48.9000 129.8000 50.2000 ;
	    RECT 130.2000 48.9000 130.6000 50.2000 ;
	    RECT 131.8000 48.9000 132.2000 50.2000 ;
	    RECT 134.2000 48.3000 134.6000 50.2000 ;
	    RECT 135.8000 48.9000 136.2000 50.2000 ;
	    RECT 138.2000 48.3000 138.6000 50.2000 ;
	    RECT 141.4000 47.9000 141.8000 50.2000 ;
	    RECT 143.8000 47.9000 144.2000 50.2000 ;
	    RECT 146.2000 48.9000 146.6000 50.2000 ;
	    RECT 1.4000 30.8000 1.8000 33.1000 ;
	    RECT 3.8000 30.8000 4.2000 33.0000 ;
	    RECT 6.6000 30.8000 7.0000 32.1000 ;
	    RECT 8.2000 30.8000 8.7000 32.1000 ;
	    RECT 11.0000 30.8000 11.4000 33.1000 ;
	    RECT 12.6000 30.8000 13.0000 32.1000 ;
	    RECT 14.2000 30.8000 14.6000 32.1000 ;
	    RECT 15.8000 30.8000 16.2000 32.1000 ;
	    RECT 16.6000 30.8000 17.0000 33.1000 ;
	    RECT 20.6000 30.8000 21.0000 33.1000 ;
	    RECT 23.8000 30.8000 24.2000 34.1000 ;
	    RECT 27.8000 30.8000 28.2000 31.9000 ;
	    RECT 29.4000 30.8000 29.8000 32.1000 ;
	    RECT 31.0000 30.8000 31.4000 32.1000 ;
	    RECT 32.6000 30.8000 33.0000 32.1000 ;
	    RECT 33.4000 30.8000 33.8000 32.1000 ;
	    RECT 35.0000 30.8000 35.4000 32.1000 ;
	    RECT 36.6000 30.8000 37.0000 32.1000 ;
	    RECT 38.2000 30.8000 38.6000 32.7000 ;
	    RECT 41.4000 30.8000 41.8000 32.9000 ;
	    RECT 43.0000 30.8000 43.4000 32.1000 ;
	    RECT 43.8000 30.8000 44.2000 33.1000 ;
	    RECT 46.2000 30.8000 46.6000 32.1000 ;
	    RECT 51.0000 30.8000 51.4000 32.7000 ;
	    RECT 54.2000 30.8000 54.6000 32.7000 ;
	    RECT 55.8000 30.8000 56.2000 32.1000 ;
	    RECT 57.4000 30.8000 57.8000 32.1000 ;
	    RECT 59.8000 30.8000 60.2000 32.7000 ;
	    RECT 61.4000 30.8000 61.8000 33.1000 ;
	    RECT 63.0000 30.8000 63.4000 33.1000 ;
	    RECT 63.8000 30.8000 64.2000 33.1000 ;
	    RECT 67.0000 30.8000 67.4000 32.1000 ;
	    RECT 68.6000 30.8000 69.0000 31.9000 ;
	    RECT 74.2000 30.8000 74.6000 33.1000 ;
	    RECT 75.0000 30.8000 75.4000 34.1000 ;
	    RECT 78.2000 30.8000 78.6000 32.1000 ;
	    RECT 80.1000 30.8000 80.5000 33.1000 ;
	    RECT 82.2000 30.8000 82.6000 32.1000 ;
	    RECT 83.0000 30.8000 83.4000 32.1000 ;
	    RECT 84.6000 30.8000 85.0000 32.1000 ;
	    RECT 87.0000 30.8000 87.4000 33.1000 ;
	    RECT 87.8000 30.8000 88.2000 32.1000 ;
	    RECT 89.4000 30.8000 89.8000 32.1000 ;
	    RECT 90.2000 30.8000 90.6000 32.1000 ;
	    RECT 91.8000 30.8000 92.2000 32.1000 ;
	    RECT 93.4000 30.8000 93.8000 32.1000 ;
	    RECT 94.2000 30.8000 94.6000 33.1000 ;
	    RECT 95.8000 30.8000 96.2000 33.1000 ;
	    RECT 99.0000 30.8000 99.4000 33.1000 ;
	    RECT 100.6000 30.8000 101.0000 33.1000 ;
	    RECT 103.0000 30.8000 103.4000 32.7000 ;
	    RECT 106.7000 30.8000 107.1000 33.0000 ;
	    RECT 109.4000 30.8000 109.8000 32.7000 ;
	    RECT 112.6000 30.8000 113.0000 33.1000 ;
	    RECT 115.3000 30.8000 115.8000 32.1000 ;
	    RECT 117.0000 30.8000 117.4000 32.1000 ;
	    RECT 119.8000 30.8000 120.2000 33.0000 ;
	    RECT 121.7000 30.8000 122.1000 33.1000 ;
	    RECT 123.8000 30.8000 124.2000 32.1000 ;
	    RECT 125.4000 30.8000 125.8000 33.1000 ;
	    RECT 128.1000 30.8000 128.6000 32.1000 ;
	    RECT 129.8000 30.8000 130.2000 32.1000 ;
	    RECT 132.6000 30.8000 133.0000 33.0000 ;
	    RECT 134.5000 30.8000 134.9000 33.1000 ;
	    RECT 136.6000 30.8000 137.0000 32.1000 ;
	    RECT 137.4000 30.8000 137.8000 32.1000 ;
	    RECT 139.0000 30.8000 139.4000 32.1000 ;
	    RECT 140.6000 30.8000 141.0000 32.1000 ;
	    RECT 142.2000 30.8000 142.6000 33.1000 ;
	    RECT 144.6000 30.8000 145.0000 33.1000 ;
	    RECT 0.2000 30.2000 148.6000 30.8000 ;
	    RECT 1.4000 28.0000 1.8000 30.2000 ;
	    RECT 4.2000 28.9000 4.6000 30.2000 ;
	    RECT 5.8000 28.9000 6.3000 30.2000 ;
	    RECT 8.6000 27.9000 9.0000 30.2000 ;
	    RECT 11.8000 28.3000 12.2000 30.2000 ;
	    RECT 15.0000 27.9000 15.4000 30.2000 ;
	    RECT 19.0000 29.1000 19.4000 30.2000 ;
	    RECT 20.6000 28.9000 21.0000 30.2000 ;
	    RECT 23.0000 28.3000 23.4000 30.2000 ;
	    RECT 25.4000 28.9000 25.8000 30.2000 ;
	    RECT 27.0000 28.9000 27.4000 30.2000 ;
	    RECT 31.0000 29.1000 31.4000 30.2000 ;
	    RECT 32.6000 28.9000 33.0000 30.2000 ;
	    RECT 34.2000 28.9000 34.6000 30.2000 ;
	    RECT 35.8000 28.9000 36.2000 30.2000 ;
	    RECT 36.9000 27.9000 37.3000 30.2000 ;
	    RECT 39.0000 28.9000 39.4000 30.2000 ;
	    RECT 40.6000 28.3000 41.0000 30.2000 ;
	    RECT 43.8000 28.9000 44.2000 30.2000 ;
	    RECT 45.4000 28.9000 45.8000 30.2000 ;
	    RECT 50.2000 28.3000 50.6000 30.2000 ;
	    RECT 51.8000 28.9000 52.2000 30.2000 ;
	    RECT 53.4000 28.9000 53.8000 30.2000 ;
	    RECT 56.6000 26.9000 57.0000 30.2000 ;
	    RECT 59.0000 28.3000 59.4000 30.2000 ;
	    RECT 60.6000 28.9000 61.0000 30.2000 ;
	    RECT 62.2000 28.9000 62.6000 30.2000 ;
	    RECT 65.4000 26.9000 65.8000 30.2000 ;
	    RECT 67.0000 28.9000 67.4000 30.2000 ;
	    RECT 68.6000 29.1000 69.0000 30.2000 ;
	    RECT 72.6000 27.9000 73.0000 30.2000 ;
	    RECT 75.8000 28.3000 76.2000 30.2000 ;
	    RECT 77.4000 28.9000 77.8000 30.2000 ;
	    RECT 79.0000 28.9000 79.4000 30.2000 ;
	    RECT 81.1000 28.0000 81.5000 30.2000 ;
	    RECT 83.8000 28.9000 84.2000 30.2000 ;
	    RECT 86.2000 27.9000 86.6000 30.2000 ;
	    RECT 87.0000 27.9000 87.4000 30.2000 ;
	    RECT 89.4000 27.9000 89.8000 30.2000 ;
	    RECT 92.1000 28.9000 92.6000 30.2000 ;
	    RECT 93.8000 28.9000 94.2000 30.2000 ;
	    RECT 96.6000 28.0000 97.0000 30.2000 ;
	    RECT 100.6000 27.9000 101.0000 30.2000 ;
	    RECT 103.0000 27.9000 103.4000 30.2000 ;
	    RECT 105.4000 28.0000 105.8000 30.2000 ;
	    RECT 108.2000 28.9000 108.6000 30.2000 ;
	    RECT 109.8000 28.9000 110.3000 30.2000 ;
	    RECT 112.6000 27.9000 113.0000 30.2000 ;
	    RECT 114.2000 28.9000 114.6000 30.2000 ;
	    RECT 115.8000 28.9000 116.2000 30.2000 ;
	    RECT 117.4000 28.9000 117.8000 30.2000 ;
	    RECT 119.0000 27.9000 119.4000 30.2000 ;
	    RECT 121.7000 28.9000 122.2000 30.2000 ;
	    RECT 123.4000 28.9000 123.8000 30.2000 ;
	    RECT 126.2000 28.0000 126.6000 30.2000 ;
	    RECT 127.8000 28.9000 128.2000 30.2000 ;
	    RECT 129.4000 28.9000 129.8000 30.2000 ;
	    RECT 130.5000 27.9000 130.9000 30.2000 ;
	    RECT 132.6000 28.9000 133.0000 30.2000 ;
	    RECT 133.4000 28.9000 133.8000 30.2000 ;
	    RECT 135.0000 28.9000 135.4000 30.2000 ;
	    RECT 136.6000 27.9000 137.0000 30.2000 ;
	    RECT 139.3000 28.9000 139.8000 30.2000 ;
	    RECT 141.0000 28.9000 141.4000 30.2000 ;
	    RECT 143.8000 28.0000 144.2000 30.2000 ;
	    RECT 146.2000 27.9000 146.6000 30.2000 ;
	    RECT 1.4000 10.8000 1.8000 13.0000 ;
	    RECT 4.2000 10.8000 4.6000 12.1000 ;
	    RECT 5.8000 10.8000 6.3000 12.1000 ;
	    RECT 8.6000 10.8000 9.0000 13.1000 ;
	    RECT 11.0000 10.8000 11.4000 13.0000 ;
	    RECT 13.8000 10.8000 14.2000 12.1000 ;
	    RECT 15.4000 10.8000 15.9000 12.1000 ;
	    RECT 18.2000 10.8000 18.6000 13.1000 ;
	    RECT 22.2000 10.8000 22.6000 14.1000 ;
	    RECT 23.8000 10.8000 24.2000 12.1000 ;
	    RECT 24.6000 10.8000 25.0000 14.1000 ;
	    RECT 27.8000 10.8000 28.2000 12.1000 ;
	    RECT 29.4000 10.8000 29.8000 12.1000 ;
	    RECT 30.2000 10.8000 30.6000 13.1000 ;
	    RECT 34.2000 10.8000 34.6000 12.7000 ;
	    RECT 35.8000 10.8000 36.2000 12.1000 ;
	    RECT 37.4000 10.8000 37.8000 12.1000 ;
	    RECT 39.0000 10.8000 39.4000 12.1000 ;
	    RECT 41.4000 10.8000 41.8000 13.1000 ;
	    RECT 42.2000 10.8000 42.6000 14.1000 ;
	    RECT 45.4000 10.8000 45.8000 12.1000 ;
	    RECT 47.0000 10.8000 47.4000 12.1000 ;
	    RECT 50.2000 10.8000 50.6000 12.7000 ;
	    RECT 55.0000 10.8000 55.4000 12.7000 ;
	    RECT 56.6000 10.8000 57.0000 13.1000 ;
	    RECT 58.5000 10.8000 58.9000 13.1000 ;
	    RECT 60.6000 10.8000 61.0000 12.1000 ;
	    RECT 61.4000 10.8000 61.8000 12.1000 ;
	    RECT 63.0000 10.8000 63.4000 12.1000 ;
	    RECT 63.8000 10.8000 64.2000 13.1000 ;
	    RECT 66.2000 10.8000 66.6000 12.1000 ;
	    RECT 67.8000 10.8000 68.2000 12.1000 ;
	    RECT 68.6000 10.8000 69.0000 12.1000 ;
	    RECT 71.8000 10.8000 72.2000 13.1000 ;
	    RECT 73.4000 10.8000 73.8000 12.1000 ;
	    RECT 75.0000 10.8000 75.4000 11.9000 ;
	    RECT 79.8000 10.8000 80.2000 12.1000 ;
	    RECT 81.4000 10.8000 81.8000 11.9000 ;
	    RECT 86.2000 10.8000 86.6000 12.1000 ;
	    RECT 87.8000 10.8000 88.2000 11.9000 ;
	    RECT 91.8000 10.8000 92.2000 12.1000 ;
	    RECT 93.4000 10.8000 93.8000 12.1000 ;
	    RECT 94.2000 10.8000 94.6000 12.1000 ;
	    RECT 95.8000 10.8000 96.2000 12.1000 ;
	    RECT 98.2000 10.8000 98.6000 13.1000 ;
	    RECT 100.9000 10.8000 101.3000 13.1000 ;
	    RECT 103.0000 10.8000 103.4000 12.1000 ;
	    RECT 103.8000 10.8000 104.2000 12.1000 ;
	    RECT 105.4000 10.8000 105.8000 12.1000 ;
	    RECT 106.2000 10.8000 106.6000 12.1000 ;
	    RECT 107.8000 10.8000 108.2000 12.1000 ;
	    RECT 108.6000 10.8000 109.0000 12.1000 ;
	    RECT 110.7000 10.8000 111.1000 13.1000 ;
	    RECT 111.8000 10.8000 112.2000 13.1000 ;
	    RECT 113.4000 10.8000 113.8000 13.1000 ;
	    RECT 115.8000 10.8000 116.2000 13.1000 ;
	    RECT 117.4000 10.8000 117.8000 13.1000 ;
	    RECT 118.2000 10.8000 118.6000 13.1000 ;
	    RECT 119.8000 10.8000 120.2000 13.1000 ;
	    RECT 121.4000 10.8000 121.8000 12.1000 ;
	    RECT 123.0000 10.8000 123.4000 12.1000 ;
	    RECT 124.6000 10.8000 125.0000 12.1000 ;
	    RECT 126.2000 10.8000 126.6000 13.0000 ;
	    RECT 129.0000 10.8000 129.4000 12.1000 ;
	    RECT 130.6000 10.8000 131.1000 12.1000 ;
	    RECT 133.4000 10.8000 133.8000 13.1000 ;
	    RECT 135.8000 10.8000 136.2000 13.1000 ;
	    RECT 138.5000 10.8000 139.0000 12.1000 ;
	    RECT 140.2000 10.8000 140.6000 12.1000 ;
	    RECT 143.0000 10.8000 143.4000 13.0000 ;
	    RECT 145.4000 10.8000 145.8000 13.1000 ;
	    RECT 147.0000 10.8000 147.4000 13.1000 ;
	    RECT 0.2000 10.2000 148.6000 10.8000 ;
	    RECT 1.4000 7.9000 1.8000 10.2000 ;
	    RECT 3.0000 7.9000 3.4000 10.2000 ;
	    RECT 4.9000 7.9000 5.3000 10.2000 ;
	    RECT 7.0000 8.9000 7.4000 10.2000 ;
	    RECT 7.8000 8.9000 8.2000 10.2000 ;
	    RECT 9.4000 8.9000 9.8000 10.2000 ;
	    RECT 11.8000 7.9000 12.2000 10.2000 ;
	    RECT 15.8000 9.1000 16.2000 10.2000 ;
	    RECT 17.4000 8.9000 17.8000 10.2000 ;
	    RECT 19.0000 8.9000 19.4000 10.2000 ;
	    RECT 20.6000 8.9000 21.0000 10.2000 ;
	    RECT 22.2000 8.9000 22.6000 10.2000 ;
	    RECT 23.8000 9.1000 24.2000 10.2000 ;
	    RECT 27.8000 7.9000 28.2000 10.2000 ;
	    RECT 30.2000 8.3000 30.6000 10.2000 ;
	    RECT 34.2000 8.3000 34.6000 10.2000 ;
	    RECT 36.6000 8.9000 37.0000 10.2000 ;
	    RECT 38.2000 9.1000 38.6000 10.2000 ;
	    RECT 42.2000 6.9000 42.6000 10.2000 ;
	    RECT 45.4000 8.9000 45.8000 10.2000 ;
	    RECT 47.0000 8.9000 47.4000 10.2000 ;
	    RECT 50.2000 8.3000 50.6000 10.2000 ;
	    RECT 53.4000 8.9000 53.8000 10.2000 ;
	    RECT 55.0000 9.1000 55.4000 10.2000 ;
	    RECT 59.8000 8.3000 60.2000 10.2000 ;
	    RECT 63.8000 7.9000 64.2000 10.2000 ;
	    RECT 65.4000 7.9000 65.8000 10.2000 ;
	    RECT 67.0000 6.9000 67.4000 10.2000 ;
	    RECT 71.0000 8.0000 71.4000 10.2000 ;
	    RECT 73.8000 8.9000 74.2000 10.2000 ;
	    RECT 75.4000 8.9000 75.9000 10.2000 ;
	    RECT 78.2000 7.9000 78.6000 10.2000 ;
	    RECT 80.6000 7.9000 81.0000 10.2000 ;
	    RECT 83.0000 7.9000 83.4000 10.2000 ;
	    RECT 85.4000 7.9000 85.8000 10.2000 ;
	    RECT 88.1000 8.9000 88.6000 10.2000 ;
	    RECT 89.8000 8.9000 90.2000 10.2000 ;
	    RECT 92.6000 8.0000 93.0000 10.2000 ;
	    RECT 95.0000 7.9000 95.4000 10.2000 ;
	    RECT 97.4000 7.9000 97.8000 10.2000 ;
	    RECT 101.4000 8.0000 101.8000 10.2000 ;
	    RECT 104.2000 8.9000 104.6000 10.2000 ;
	    RECT 105.8000 8.9000 106.3000 10.2000 ;
	    RECT 108.6000 7.9000 109.0000 10.2000 ;
	    RECT 111.0000 7.9000 111.4000 10.2000 ;
	    RECT 113.4000 7.9000 113.8000 10.2000 ;
	    RECT 115.8000 7.9000 116.2000 10.2000 ;
	    RECT 118.2000 7.9000 118.6000 10.2000 ;
	    RECT 120.6000 7.9000 121.0000 10.2000 ;
	    RECT 123.0000 7.9000 123.4000 10.2000 ;
	    RECT 125.4000 7.9000 125.8000 10.2000 ;
	    RECT 127.9000 9.9000 128.3000 10.2000 ;
	    RECT 127.8000 8.2000 128.3000 9.9000 ;
	    RECT 130.9000 8.2000 131.4000 10.2000 ;
	    RECT 133.4000 7.9000 133.8000 10.2000 ;
	    RECT 135.8000 7.9000 136.2000 10.2000 ;
	    RECT 138.2000 7.9000 138.6000 10.2000 ;
	    RECT 140.6000 7.9000 141.0000 10.2000 ;
	    RECT 143.0000 7.9000 143.4000 10.2000 ;
	    RECT 144.6000 7.9000 145.0000 10.2000 ;
         LAYER metal2 ;
	    RECT 97.6000 110.3000 99.2000 110.7000 ;
	    RECT 97.6000 90.3000 99.2000 90.7000 ;
	    RECT 97.6000 70.3000 99.2000 70.7000 ;
	    RECT 97.6000 50.3000 99.2000 50.7000 ;
	    RECT 97.6000 30.3000 99.2000 30.7000 ;
	    RECT 97.6000 10.3000 99.2000 10.7000 ;
         LAYER metal3 ;
	    RECT 97.6000 110.3000 99.2000 110.7000 ;
	    RECT 97.6000 90.3000 99.2000 90.7000 ;
	    RECT 97.6000 70.3000 99.2000 70.7000 ;
	    RECT 97.6000 50.3000 99.2000 50.7000 ;
	    RECT 97.6000 30.3000 99.2000 30.7000 ;
	    RECT 97.6000 10.3000 99.2000 10.7000 ;
         LAYER metal4 ;
	    RECT 97.6000 110.3000 99.2000 110.7000 ;
	    RECT 97.6000 90.3000 99.2000 90.7000 ;
	    RECT 97.6000 70.3000 99.2000 70.7000 ;
	    RECT 97.6000 50.3000 99.2000 50.7000 ;
	    RECT 97.6000 30.3000 99.2000 30.7000 ;
	    RECT 97.6000 10.3000 99.2000 10.7000 ;
         LAYER metal5 ;
	    RECT 97.6000 110.2000 99.2000 110.7000 ;
	    RECT 97.6000 90.2000 99.2000 90.7000 ;
	    RECT 97.6000 70.2000 99.2000 70.7000 ;
	    RECT 97.6000 50.2000 99.2000 50.7000 ;
	    RECT 97.6000 30.2000 99.2000 30.7000 ;
	    RECT 97.6000 10.2000 99.2000 10.7000 ;
         LAYER metal6 ;
	    RECT 97.6000 -3.0000 99.2000 123.0000 ;
      END
   END gnd
   PIN clk
      PORT
         LAYER metal1 ;
	    RECT 21.5000 86.2000 21.9000 86.6000 ;
	    RECT 93.5000 86.2000 93.9000 86.6000 ;
	    RECT 101.5000 86.2000 101.9000 86.6000 ;
	    RECT 21.4000 85.8000 21.9000 86.2000 ;
	    RECT 93.4000 85.8000 93.9000 86.2000 ;
	    RECT 101.4000 85.8000 101.9000 86.2000 ;
	    RECT 19.7000 46.2000 20.1000 46.6000 ;
	    RECT 19.7000 45.8000 20.2000 46.2000 ;
	    RECT 96.5000 35.1000 97.0000 35.2000 ;
	    RECT 98.2000 35.1000 98.6000 35.2000 ;
	    RECT 96.5000 34.8000 98.6000 35.1000 ;
	    RECT 101.3000 34.8000 101.8000 35.2000 ;
	    RECT 96.5000 34.4000 96.9000 34.8000 ;
	    RECT 101.3000 34.4000 101.7000 34.8000 ;
         LAYER metal2 ;
	    RECT 21.4000 86.1000 21.8000 86.2000 ;
	    RECT 93.4000 86.1000 93.8000 86.2000 ;
	    RECT 94.2000 86.1000 94.6000 86.2000 ;
	    RECT 21.4000 85.8000 22.5000 86.1000 ;
	    RECT 93.4000 85.8000 94.6000 86.1000 ;
	    RECT 101.4000 85.8000 101.8000 86.2000 ;
	    RECT 22.2000 82.2000 22.5000 85.8000 ;
	    RECT 94.2000 82.2000 94.5000 85.8000 ;
	    RECT 22.2000 81.8000 22.6000 82.2000 ;
	    RECT 94.2000 81.8000 94.6000 82.2000 ;
	    RECT 101.4000 74.2000 101.7000 85.8000 ;
	    RECT 101.4000 73.8000 101.8000 74.2000 ;
	    RECT 19.8000 46.8000 20.2000 47.2000 ;
	    RECT 19.8000 46.2000 20.1000 46.8000 ;
	    RECT 19.8000 45.8000 20.2000 46.2000 ;
	    RECT 98.2000 35.1000 98.6000 35.2000 ;
	    RECT 99.0000 35.1000 99.4000 35.2000 ;
	    RECT 98.2000 34.8000 99.4000 35.1000 ;
	    RECT 100.6000 35.1000 101.0000 35.2000 ;
	    RECT 101.4000 35.1000 101.8000 35.2000 ;
	    RECT 100.6000 34.8000 101.8000 35.1000 ;
         LAYER metal3 ;
	    RECT 94.2000 86.1000 94.6000 86.2000 ;
	    RECT 101.4000 86.1000 101.8000 86.2000 ;
	    RECT 94.2000 85.8000 101.8000 86.1000 ;
	    RECT 19.8000 82.1000 20.2000 82.2000 ;
	    RECT 22.2000 82.1000 22.6000 82.2000 ;
	    RECT 94.2000 82.1000 94.6000 82.2000 ;
	    RECT 19.8000 81.8000 94.6000 82.1000 ;
	    RECT 100.6000 74.1000 101.0000 74.2000 ;
	    RECT 101.4000 74.1000 101.8000 74.2000 ;
	    RECT 100.6000 73.8000 101.8000 74.1000 ;
	    RECT 19.8000 46.8000 20.2000 47.2000 ;
	    RECT 19.8000 46.1000 20.1000 46.8000 ;
	    RECT 20.6000 46.1000 21.0000 46.2000 ;
	    RECT -2.6000 45.8000 21.0000 46.1000 ;
	    RECT 99.0000 35.1000 99.4000 35.2000 ;
	    RECT 100.6000 35.1000 101.0000 35.2000 ;
	    RECT 99.0000 34.8000 101.0000 35.1000 ;
         LAYER metal4 ;
	    RECT 19.8000 81.8000 20.2000 82.2000 ;
	    RECT 19.8000 46.1000 20.1000 81.8000 ;
	    RECT 100.6000 73.8000 101.0000 74.2000 ;
	    RECT 20.6000 46.1000 21.0000 46.2000 ;
	    RECT 19.8000 45.8000 21.0000 46.1000 ;
	    RECT 100.6000 35.2000 100.9000 73.8000 ;
	    RECT 100.6000 34.8000 101.0000 35.2000 ;
      END
   END clk
   PIN INPD<0>
      PORT
         LAYER metal1 ;
	    RECT 92.6000 46.8000 93.0000 47.2000 ;
	    RECT 92.6000 46.6000 92.9000 46.8000 ;
	    RECT 92.5000 46.2000 92.9000 46.6000 ;
         LAYER metal2 ;
	    RECT 92.6000 46.8000 93.0000 47.2000 ;
	    RECT 92.6000 45.1000 92.9000 46.8000 ;
	    RECT 93.4000 45.1000 93.8000 45.2000 ;
	    RECT 92.6000 44.8000 93.8000 45.1000 ;
	    RECT 91.8000 0.8000 92.2000 1.2000 ;
	    RECT 91.8000 -2.2000 92.1000 0.8000 ;
         LAYER metal3 ;
	    RECT 92.6000 45.1000 93.0000 45.2000 ;
	    RECT 93.4000 45.1000 93.8000 45.2000 ;
	    RECT 92.6000 44.8000 93.8000 45.1000 ;
	    RECT 91.8000 1.1000 92.2000 1.2000 ;
	    RECT 92.6000 1.1000 93.0000 1.2000 ;
	    RECT 91.8000 0.8000 93.0000 1.1000 ;
         LAYER metal4 ;
	    RECT 92.6000 44.8000 93.0000 45.2000 ;
	    RECT 92.6000 1.2000 92.9000 44.8000 ;
	    RECT 92.6000 0.8000 93.0000 1.2000 ;
      END
   END INPD<0>
   PIN INPD<1>
      PORT
         LAYER metal1 ;
	    RECT 110.2000 105.8000 110.6000 106.6000 ;
         LAYER metal2 ;
	    RECT 111.8000 120.2000 112.1000 123.1000 ;
	    RECT 110.2000 119.8000 110.6000 120.2000 ;
	    RECT 111.8000 119.8000 112.2000 120.2000 ;
	    RECT 110.2000 106.2000 110.5000 119.8000 ;
	    RECT 110.2000 105.8000 110.6000 106.2000 ;
         LAYER metal3 ;
	    RECT 110.2000 120.1000 110.6000 120.2000 ;
	    RECT 111.8000 120.1000 112.2000 120.2000 ;
	    RECT 110.2000 119.8000 112.2000 120.1000 ;
      END
   END INPD<1>
   PIN INPD<2>
      PORT
         LAYER metal1 ;
	    RECT 118.2000 105.8000 118.6000 106.6000 ;
         LAYER metal2 ;
	    RECT 118.2000 122.8000 119.3000 123.1000 ;
	    RECT 119.0000 111.1000 119.3000 122.8000 ;
	    RECT 118.2000 110.8000 119.3000 111.1000 ;
	    RECT 118.2000 106.2000 118.5000 110.8000 ;
	    RECT 118.2000 105.8000 118.6000 106.2000 ;
      END
   END INPD<2>
   PIN INPD<3>
      PORT
         LAYER metal1 ;
	    RECT 144.6000 67.8000 145.0000 68.6000 ;
         LAYER metal2 ;
	    RECT 144.6000 77.8000 145.0000 78.2000 ;
	    RECT 144.6000 68.2000 144.9000 77.8000 ;
	    RECT 144.6000 67.8000 145.0000 68.2000 ;
         LAYER metal3 ;
	    RECT 144.6000 78.1000 145.0000 78.2000 ;
	    RECT 144.6000 77.8000 151.3000 78.1000 ;
      END
   END INPD<3>
   PIN INPD<4>
      PORT
         LAYER metal1 ;
	    RECT 140.6000 67.8000 141.0000 68.6000 ;
         LAYER metal2 ;
	    RECT 141.4000 75.8000 141.8000 76.2000 ;
	    RECT 141.4000 72.1000 141.7000 75.8000 ;
	    RECT 140.6000 71.8000 141.7000 72.1000 ;
	    RECT 140.6000 68.2000 140.9000 71.8000 ;
	    RECT 140.6000 67.8000 141.0000 68.2000 ;
         LAYER metal3 ;
	    RECT 141.4000 76.1000 141.8000 76.2000 ;
	    RECT 141.4000 75.8000 151.3000 76.1000 ;
      END
   END INPD<4>
   PIN INPD<5>
      PORT
         LAYER metal1 ;
	    RECT 146.2000 48.1000 146.6000 48.6000 ;
	    RECT 147.0000 48.1000 147.4000 48.2000 ;
	    RECT 146.2000 47.8000 147.4000 48.1000 ;
         LAYER metal2 ;
	    RECT 147.0000 71.8000 147.4000 72.2000 ;
	    RECT 147.0000 48.2000 147.3000 71.8000 ;
	    RECT 147.0000 47.8000 147.4000 48.2000 ;
         LAYER metal3 ;
	    RECT 147.0000 72.1000 147.4000 72.2000 ;
	    RECT 147.0000 71.8000 151.3000 72.1000 ;
      END
   END INPD<5>
   PIN INPD<6>
      PORT
         LAYER metal1 ;
	    RECT 143.8000 92.4000 144.2000 93.2000 ;
         LAYER metal2 ;
	    RECT 143.8000 95.8000 144.2000 96.2000 ;
	    RECT 143.8000 93.2000 144.1000 95.8000 ;
	    RECT 143.8000 92.8000 144.2000 93.2000 ;
         LAYER metal3 ;
	    RECT 143.8000 96.1000 144.2000 96.2000 ;
	    RECT 143.8000 95.8000 151.3000 96.1000 ;
      END
   END INPD<6>
   PIN INPD<7>
      PORT
         LAYER metal1 ;
	    RECT 137.4000 52.4000 137.8000 53.2000 ;
         LAYER metal2 ;
	    RECT 137.4000 52.8000 137.8000 53.2000 ;
	    RECT 137.4000 52.2000 137.7000 52.8000 ;
	    RECT 137.4000 51.8000 137.8000 52.2000 ;
         LAYER metal3 ;
	    RECT 137.4000 52.1000 137.8000 52.2000 ;
	    RECT 151.0000 52.1000 151.3000 53.1000 ;
	    RECT 137.4000 51.8000 151.3000 52.1000 ;
      END
   END INPD<7>
   PIN INPD<8>
   END INPD<8>
   PIN INPD<9>
   END INPD<9>
   PIN INPD<10>
   END INPD<10>
   PIN INPD<11>
   END INPD<11>
   PIN INPD<12>
   END INPD<12>
   PIN INPD<13>
   END INPD<13>
   PIN INPD<14>
   END INPD<14>
   PIN INPD<15>
   END INPD<15>
   PIN RDATA<0>
      PORT
         LAYER metal1 ;
	    RECT 88.6000 45.8000 89.0000 46.6000 ;
         LAYER metal2 ;
	    RECT 87.8000 47.1000 88.2000 47.2000 ;
	    RECT 87.8000 46.8000 88.9000 47.1000 ;
	    RECT 88.6000 46.2000 88.9000 46.8000 ;
	    RECT 88.6000 45.8000 89.0000 46.2000 ;
	    RECT 88.6000 0.8000 89.0000 1.2000 ;
	    RECT 88.6000 -2.2000 88.9000 0.8000 ;
         LAYER metal3 ;
	    RECT 87.8000 47.1000 88.2000 47.2000 ;
	    RECT 88.6000 47.1000 89.0000 47.2000 ;
	    RECT 87.8000 46.8000 89.0000 47.1000 ;
	    RECT 88.6000 1.8000 89.0000 2.2000 ;
	    RECT 88.6000 1.2000 88.9000 1.8000 ;
	    RECT 88.6000 0.8000 89.0000 1.2000 ;
         LAYER metal4 ;
	    RECT 88.6000 46.8000 89.0000 47.2000 ;
	    RECT 88.6000 2.2000 88.9000 46.8000 ;
	    RECT 88.6000 1.8000 89.0000 2.2000 ;
      END
   END RDATA<0>
   PIN RDATA<1>
      PORT
         LAYER metal1 ;
	    RECT 109.4000 117.1000 109.8000 117.2000 ;
	    RECT 108.6000 116.8000 109.8000 117.1000 ;
	    RECT 108.6000 115.8000 109.0000 116.8000 ;
         LAYER metal2 ;
	    RECT 109.4000 117.2000 109.7000 123.1000 ;
	    RECT 109.4000 116.8000 109.8000 117.2000 ;
      END
   END RDATA<1>
   PIN RDATA<2>
      PORT
         LAYER metal1 ;
	    RECT 147.8000 57.1000 148.2000 57.2000 ;
	    RECT 147.0000 56.8000 148.2000 57.1000 ;
	    RECT 147.0000 55.8000 147.4000 56.8000 ;
         LAYER metal2 ;
	    RECT 147.8000 73.8000 148.2000 74.2000 ;
	    RECT 147.8000 57.2000 148.1000 73.8000 ;
	    RECT 147.8000 56.8000 148.2000 57.2000 ;
         LAYER metal3 ;
	    RECT 147.8000 74.1000 148.2000 74.2000 ;
	    RECT 147.8000 73.8000 151.3000 74.1000 ;
      END
   END RDATA<2>
   PIN RDATA<3>
      PORT
         LAYER metal1 ;
	    RECT 142.2000 55.8000 142.6000 57.2000 ;
         LAYER metal2 ;
	    RECT 142.2000 59.8000 142.6000 60.2000 ;
	    RECT 142.2000 57.2000 142.5000 59.8000 ;
	    RECT 142.2000 56.8000 142.6000 57.2000 ;
         LAYER metal3 ;
	    RECT 142.2000 60.1000 142.6000 60.2000 ;
	    RECT 142.2000 59.8000 151.3000 60.1000 ;
      END
   END RDATA<3>
   PIN RDATA<4>
      PORT
         LAYER metal1 ;
	    RECT 129.4000 55.8000 129.8000 57.2000 ;
         LAYER metal2 ;
	    RECT 129.4000 63.8000 129.8000 64.2000 ;
	    RECT 129.4000 57.2000 129.7000 63.8000 ;
	    RECT 129.4000 56.8000 129.8000 57.2000 ;
         LAYER metal3 ;
	    RECT 148.6000 66.1000 149.0000 66.2000 ;
	    RECT 148.6000 65.8000 151.3000 66.1000 ;
	    RECT 129.4000 64.1000 129.8000 64.2000 ;
	    RECT 148.6000 64.1000 149.0000 64.2000 ;
	    RECT 129.4000 63.8000 149.0000 64.1000 ;
         LAYER metal4 ;
	    RECT 148.6000 65.8000 149.0000 66.2000 ;
	    RECT 148.6000 64.2000 148.9000 65.8000 ;
	    RECT 148.6000 63.8000 149.0000 64.2000 ;
      END
   END RDATA<4>
   PIN RDATA<5>
      PORT
         LAYER metal1 ;
	    RECT 146.2000 5.1000 146.6000 5.2000 ;
	    RECT 148.6000 5.1000 149.0000 5.2000 ;
	    RECT 146.2000 4.8000 149.0000 5.1000 ;
	    RECT 146.2000 4.4000 146.6000 4.8000 ;
         LAYER metal2 ;
	    RECT 148.6000 15.8000 149.0000 16.2000 ;
	    RECT 148.6000 5.2000 148.9000 15.8000 ;
	    RECT 148.6000 4.8000 149.0000 5.2000 ;
         LAYER metal3 ;
	    RECT 148.6000 16.1000 149.0000 16.2000 ;
	    RECT 148.6000 15.8000 151.3000 16.1000 ;
      END
   END RDATA<5>
   PIN RDATA<6>
      PORT
         LAYER metal1 ;
	    RECT 111.0000 115.8000 111.4000 117.2000 ;
         LAYER metal2 ;
	    RECT 113.4000 119.2000 113.7000 123.1000 ;
	    RECT 111.0000 118.8000 111.4000 119.2000 ;
	    RECT 113.4000 118.8000 113.8000 119.2000 ;
	    RECT 111.0000 117.2000 111.3000 118.8000 ;
	    RECT 111.0000 116.8000 111.4000 117.2000 ;
         LAYER metal3 ;
	    RECT 111.0000 119.1000 111.4000 119.2000 ;
	    RECT 113.4000 119.1000 113.8000 119.2000 ;
	    RECT 111.0000 118.8000 113.8000 119.1000 ;
      END
   END RDATA<6>
   PIN RDATA<7>
      PORT
         LAYER metal1 ;
	    RECT 143.0000 64.4000 143.4000 65.2000 ;
         LAYER metal2 ;
	    RECT 143.0000 67.8000 143.4000 68.2000 ;
	    RECT 143.0000 65.2000 143.3000 67.8000 ;
	    RECT 143.0000 64.8000 143.4000 65.2000 ;
         LAYER metal3 ;
	    RECT 143.0000 68.1000 143.4000 68.2000 ;
	    RECT 143.0000 67.8000 151.3000 68.1000 ;
      END
   END RDATA<7>
   PIN RF
      PORT
         LAYER metal1 ;
	    RECT 42.2000 4.8000 42.6000 5.6000 ;
         LAYER metal2 ;
	    RECT 42.2000 4.8000 42.6000 5.2000 ;
	    RECT 42.2000 -2.2000 42.5000 4.8000 ;
      END
   END RF
   PIN WF
      PORT
         LAYER metal1 ;
	    RECT 3.0000 6.8000 3.4000 7.6000 ;
         LAYER metal2 ;
	    RECT 3.0000 7.8000 3.4000 8.2000 ;
	    RECT 3.0000 7.2000 3.3000 7.8000 ;
	    RECT 3.0000 6.8000 3.4000 7.2000 ;
         LAYER metal3 ;
	    RECT 3.0000 8.1000 3.4000 8.2000 ;
	    RECT -2.6000 7.8000 3.4000 8.1000 ;
      END
   END WF
   PIN NEXTOP<0>
      PORT
         LAYER metal1 ;
	    RECT 43.8000 33.4000 44.2000 34.2000 ;
	    RECT 36.6000 32.4000 37.0000 33.2000 ;
	    RECT 55.8000 32.4000 56.2000 33.2000 ;
	    RECT 23.0000 25.8000 23.4000 26.6000 ;
	    RECT 42.2000 17.1000 42.6000 17.2000 ;
	    RECT 43.0000 17.1000 43.4000 17.2000 ;
	    RECT 43.8000 17.1000 44.2000 17.2000 ;
	    RECT 42.2000 16.8000 44.2000 17.1000 ;
	    RECT 43.8000 16.4000 44.2000 16.8000 ;
	    RECT 23.8000 16.1000 24.2000 16.2000 ;
	    RECT 24.6000 16.1000 25.0000 16.2000 ;
	    RECT 23.8000 15.8000 25.0000 16.1000 ;
	    RECT 24.6000 15.4000 25.0000 15.8000 ;
	    RECT 55.0000 15.1000 55.4000 15.2000 ;
	    RECT 55.8000 15.1000 56.2000 15.2000 ;
	    RECT 55.0000 14.8000 56.2000 15.1000 ;
	    RECT 55.0000 14.4000 55.4000 14.8000 ;
	    RECT 20.6000 7.8000 21.0000 8.6000 ;
	    RECT 36.6000 7.8000 37.5000 8.2000 ;
         LAYER metal2 ;
	    RECT 36.6000 33.8000 37.0000 34.2000 ;
	    RECT 43.8000 33.8000 44.2000 34.2000 ;
	    RECT 55.8000 33.8000 56.2000 34.2000 ;
	    RECT 36.6000 33.2000 36.9000 33.8000 ;
	    RECT 43.8000 33.2000 44.1000 33.8000 ;
	    RECT 55.8000 33.2000 56.1000 33.8000 ;
	    RECT 36.6000 32.8000 37.0000 33.2000 ;
	    RECT 43.8000 32.8000 44.2000 33.2000 ;
	    RECT 55.8000 32.8000 56.2000 33.2000 ;
	    RECT 43.8000 31.1000 44.1000 32.8000 ;
	    RECT 43.0000 30.8000 44.1000 31.1000 ;
	    RECT 23.0000 25.8000 23.4000 26.2000 ;
	    RECT 23.0000 22.1000 23.3000 25.8000 ;
	    RECT 23.0000 21.8000 24.1000 22.1000 ;
	    RECT 23.8000 16.2000 24.1000 21.8000 ;
	    RECT 43.0000 17.2000 43.3000 30.8000 ;
	    RECT 42.2000 16.8000 42.6000 17.2000 ;
	    RECT 43.0000 16.8000 43.4000 17.2000 ;
	    RECT 55.8000 16.8000 56.2000 17.2000 ;
	    RECT 23.8000 15.8000 24.2000 16.2000 ;
	    RECT 23.8000 14.2000 24.1000 15.8000 ;
	    RECT 20.6000 13.8000 21.0000 14.2000 ;
	    RECT 23.8000 13.8000 24.2000 14.2000 ;
	    RECT 20.6000 8.2000 20.9000 13.8000 ;
	    RECT 42.2000 8.2000 42.5000 16.8000 ;
	    RECT 55.8000 15.2000 56.1000 16.8000 ;
	    RECT 55.8000 14.8000 56.2000 15.2000 ;
	    RECT 20.6000 7.8000 21.0000 8.2000 ;
	    RECT 35.8000 8.1000 36.2000 8.2000 ;
	    RECT 36.6000 8.1000 37.0000 8.2000 ;
	    RECT 35.8000 7.8000 37.0000 8.1000 ;
	    RECT 42.2000 7.8000 42.6000 8.2000 ;
	    RECT 36.6000 -2.2000 36.9000 7.8000 ;
         LAYER metal3 ;
	    RECT 36.6000 33.8000 37.0000 34.2000 ;
	    RECT 43.8000 34.1000 44.2000 34.2000 ;
	    RECT 55.8000 34.1000 56.2000 34.2000 ;
	    RECT 43.8000 33.8000 56.2000 34.1000 ;
	    RECT 36.6000 33.1000 36.9000 33.8000 ;
	    RECT 43.8000 33.1000 44.2000 33.2000 ;
	    RECT 36.6000 32.8000 44.2000 33.1000 ;
	    RECT 42.2000 17.1000 42.6000 17.2000 ;
	    RECT 55.8000 17.1000 56.2000 17.2000 ;
	    RECT 42.2000 16.8000 56.2000 17.1000 ;
	    RECT 20.6000 14.1000 21.0000 14.2000 ;
	    RECT 23.8000 14.1000 24.2000 14.2000 ;
	    RECT 20.6000 13.8000 24.2000 14.1000 ;
	    RECT 20.6000 8.1000 21.0000 8.2000 ;
	    RECT 35.8000 8.1000 36.2000 8.2000 ;
	    RECT 42.2000 8.1000 42.6000 8.2000 ;
	    RECT 20.6000 7.8000 42.6000 8.1000 ;
      END
   END NEXTOP<0>
   PIN NEXTOP<1>
      PORT
         LAYER metal1 ;
	    RECT 38.9000 28.2000 39.3000 28.6000 ;
	    RECT 39.0000 27.8000 39.4000 28.2000 ;
	    RECT 57.4000 25.1000 57.8000 25.2000 ;
	    RECT 57.4000 24.8000 58.1000 25.1000 ;
	    RECT 57.8000 24.2000 58.1000 24.8000 ;
	    RECT 56.6000 24.1000 57.0000 24.2000 ;
	    RECT 57.8000 24.1000 58.2000 24.2000 ;
	    RECT 56.6000 23.8000 58.2000 24.1000 ;
	    RECT 39.0000 16.1000 39.4000 16.2000 ;
	    RECT 39.8000 16.1000 40.2000 16.6000 ;
	    RECT 39.0000 15.8000 40.2000 16.1000 ;
	    RECT 43.0000 14.8000 43.8000 15.2000 ;
	    RECT 45.4000 14.8000 45.8000 15.6000 ;
	    RECT 56.6000 13.4000 57.0000 14.2000 ;
	    RECT 71.8000 13.4000 72.2000 14.2000 ;
         LAYER metal2 ;
	    RECT 39.0000 28.8000 39.4000 29.2000 ;
	    RECT 39.0000 28.2000 39.3000 28.8000 ;
	    RECT 39.0000 27.8000 39.4000 28.2000 ;
	    RECT 56.6000 23.8000 57.0000 24.2000 ;
	    RECT 39.0000 16.1000 39.4000 16.2000 ;
	    RECT 39.8000 16.1000 40.2000 16.2000 ;
	    RECT 39.0000 15.8000 40.2000 16.1000 ;
	    RECT 43.0000 15.8000 43.4000 16.2000 ;
	    RECT 45.4000 15.8000 45.8000 16.2000 ;
	    RECT 47.8000 15.8000 48.2000 16.2000 ;
	    RECT 43.0000 15.2000 43.3000 15.8000 ;
	    RECT 45.4000 15.2000 45.7000 15.8000 ;
	    RECT 43.0000 14.8000 43.4000 15.2000 ;
	    RECT 45.4000 14.8000 45.8000 15.2000 ;
	    RECT 47.8000 10.2000 48.1000 15.8000 ;
	    RECT 56.6000 14.2000 56.9000 23.8000 ;
	    RECT 56.6000 13.8000 57.0000 14.2000 ;
	    RECT 71.8000 13.8000 72.2000 14.2000 ;
	    RECT 56.6000 10.2000 56.9000 13.8000 ;
	    RECT 71.8000 10.2000 72.1000 13.8000 ;
	    RECT 47.8000 9.8000 48.2000 10.2000 ;
	    RECT 56.6000 9.8000 57.0000 10.2000 ;
	    RECT 71.8000 9.8000 72.2000 10.2000 ;
	    RECT 71.8000 -2.2000 72.1000 9.8000 ;
         LAYER metal3 ;
	    RECT 39.0000 29.1000 39.4000 29.2000 ;
	    RECT 39.8000 29.1000 40.2000 29.2000 ;
	    RECT 39.0000 28.8000 40.2000 29.1000 ;
	    RECT 39.0000 16.1000 39.4000 16.2000 ;
	    RECT 39.8000 16.1000 40.2000 16.2000 ;
	    RECT 43.0000 16.1000 43.4000 16.2000 ;
	    RECT 45.4000 16.1000 45.8000 16.2000 ;
	    RECT 47.8000 16.1000 48.2000 16.2000 ;
	    RECT 39.0000 15.8000 48.2000 16.1000 ;
	    RECT 47.8000 10.1000 48.2000 10.2000 ;
	    RECT 56.6000 10.1000 57.0000 10.2000 ;
	    RECT 71.8000 10.1000 72.2000 10.2000 ;
	    RECT 47.8000 9.8000 72.2000 10.1000 ;
         LAYER metal4 ;
	    RECT 39.8000 29.1000 40.2000 29.2000 ;
	    RECT 39.0000 28.8000 40.2000 29.1000 ;
	    RECT 39.0000 16.2000 39.3000 28.8000 ;
	    RECT 39.0000 15.8000 39.4000 16.2000 ;
      END
   END NEXTOP<1>
   PIN NEXTOP<2>
      PORT
         LAYER metal1 ;
	    RECT 62.2000 27.8000 62.6000 28.6000 ;
	    RECT 36.6000 26.1000 37.0000 26.2000 ;
	    RECT 36.6000 25.8000 37.4000 26.1000 ;
	    RECT 37.0000 25.6000 37.4000 25.8000 ;
	    RECT 41.4000 16.1000 41.8000 16.2000 ;
	    RECT 42.2000 16.1000 42.6000 16.2000 ;
	    RECT 41.4000 15.8000 42.6000 16.1000 ;
	    RECT 42.2000 15.4000 42.6000 15.8000 ;
	    RECT 41.4000 13.4000 41.8000 14.2000 ;
	    RECT 47.0000 12.4000 47.4000 13.2000 ;
	    RECT 67.8000 13.1000 68.2000 13.2000 ;
	    RECT 68.6000 13.1000 69.0000 13.2000 ;
	    RECT 67.8000 12.8000 69.0000 13.1000 ;
	    RECT 67.8000 12.4000 68.2000 12.8000 ;
	    RECT 68.6000 12.4000 69.0000 12.8000 ;
	    RECT 61.4000 5.1000 61.8000 5.2000 ;
	    RECT 61.1000 4.8000 61.8000 5.1000 ;
	    RECT 61.1000 4.2000 61.4000 4.8000 ;
	    RECT 61.0000 3.8000 61.4000 4.2000 ;
         LAYER metal2 ;
	    RECT 62.2000 27.8000 62.6000 28.2000 ;
	    RECT 36.6000 25.8000 37.0000 26.2000 ;
	    RECT 36.6000 14.2000 36.9000 25.8000 ;
	    RECT 41.4000 15.8000 41.8000 16.2000 ;
	    RECT 41.4000 14.2000 41.7000 15.8000 ;
	    RECT 62.2000 14.2000 62.5000 27.8000 ;
	    RECT 36.6000 13.8000 37.0000 14.2000 ;
	    RECT 41.4000 13.8000 41.8000 14.2000 ;
	    RECT 47.0000 13.8000 47.4000 14.2000 ;
	    RECT 61.4000 13.8000 61.8000 14.2000 ;
	    RECT 62.2000 13.8000 62.6000 14.2000 ;
	    RECT 67.8000 13.8000 68.2000 14.2000 ;
	    RECT 47.0000 13.2000 47.3000 13.8000 ;
	    RECT 47.0000 12.8000 47.4000 13.2000 ;
	    RECT 61.4000 5.2000 61.7000 13.8000 ;
	    RECT 67.8000 13.2000 68.1000 13.8000 ;
	    RECT 67.8000 12.8000 68.2000 13.2000 ;
	    RECT 61.4000 4.8000 61.8000 5.2000 ;
	    RECT 61.4000 -2.2000 61.7000 4.8000 ;
         LAYER metal3 ;
	    RECT 36.6000 14.1000 37.0000 14.2000 ;
	    RECT 41.4000 14.1000 41.8000 14.2000 ;
	    RECT 47.0000 14.1000 47.4000 14.2000 ;
	    RECT 61.4000 14.1000 61.8000 14.2000 ;
	    RECT 62.2000 14.1000 62.6000 14.2000 ;
	    RECT 67.8000 14.1000 68.2000 14.2000 ;
	    RECT 36.6000 13.8000 68.2000 14.1000 ;
      END
   END NEXTOP<2>
   PIN IR
      PORT
         LAYER metal1 ;
	    RECT 103.8000 115.9000 104.2000 119.9000 ;
	    RECT 103.9000 114.8000 104.2000 115.9000 ;
	    RECT 103.8000 111.1000 104.2000 114.8000 ;
         LAYER metal2 ;
	    RECT 105.4000 121.2000 105.7000 123.1000 ;
	    RECT 103.8000 120.8000 104.2000 121.2000 ;
	    RECT 105.4000 120.8000 105.8000 121.2000 ;
	    RECT 103.8000 119.2000 104.1000 120.8000 ;
	    RECT 103.8000 118.8000 104.2000 119.2000 ;
         LAYER metal3 ;
	    RECT 103.8000 121.1000 104.2000 121.2000 ;
	    RECT 105.4000 121.1000 105.8000 121.2000 ;
	    RECT 103.8000 120.8000 105.8000 121.1000 ;
      END
   END IR
   PIN OW
      PORT
         LAYER metal1 ;
	    RECT 134.2000 6.2000 134.6000 9.9000 ;
	    RECT 134.3000 5.1000 134.6000 6.2000 ;
	    RECT 134.2000 1.1000 134.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 134.2000 1.8000 134.6000 2.2000 ;
	    RECT 134.2000 -2.2000 134.5000 1.8000 ;
      END
   END OW
   PIN OUTPD<0>
      PORT
         LAYER metal1 ;
	    RECT 95.8000 6.2000 96.2000 9.9000 ;
	    RECT 95.9000 5.1000 96.2000 6.2000 ;
	    RECT 95.8000 1.1000 96.2000 5.1000 ;
         LAYER metal2 ;
	    RECT 95.8000 1.8000 96.2000 2.2000 ;
	    RECT 95.8000 -2.2000 96.1000 1.8000 ;
      END
   END OUTPD<0>
   PIN OUTPD<1>
      PORT
         LAYER metal1 ;
	    RECT 123.0000 115.9000 123.4000 119.9000 ;
	    RECT 123.1000 114.8000 123.4000 115.9000 ;
	    RECT 123.0000 111.1000 123.4000 114.8000 ;
         LAYER metal2 ;
	    RECT 123.0000 119.2000 123.3000 123.1000 ;
	    RECT 123.0000 118.8000 123.4000 119.2000 ;
      END
   END OUTPD<1>
   PIN OUTPD<2>
      PORT
         LAYER metal1 ;
	    RECT 123.8000 115.9000 124.2000 119.9000 ;
	    RECT 123.8000 114.8000 124.1000 115.9000 ;
	    RECT 123.8000 111.1000 124.2000 114.8000 ;
         LAYER metal2 ;
	    RECT 125.4000 121.2000 125.7000 123.1000 ;
	    RECT 123.8000 120.8000 124.2000 121.2000 ;
	    RECT 125.4000 120.8000 125.8000 121.2000 ;
	    RECT 123.8000 119.2000 124.1000 120.8000 ;
	    RECT 123.8000 118.8000 124.2000 119.2000 ;
         LAYER metal3 ;
	    RECT 123.8000 121.1000 124.2000 121.2000 ;
	    RECT 125.4000 121.1000 125.8000 121.2000 ;
	    RECT 123.8000 120.8000 125.8000 121.1000 ;
      END
   END OUTPD<2>
   PIN OUTPD<3>
      PORT
         LAYER metal1 ;
	    RECT 143.0000 35.9000 143.4000 39.9000 ;
	    RECT 143.1000 34.8000 143.4000 35.9000 ;
	    RECT 143.0000 31.1000 143.4000 34.8000 ;
         LAYER metal2 ;
	    RECT 143.0000 38.8000 143.4000 39.2000 ;
	    RECT 143.0000 38.2000 143.3000 38.8000 ;
	    RECT 143.0000 37.8000 143.4000 38.2000 ;
         LAYER metal3 ;
	    RECT 143.0000 38.8000 143.4000 39.2000 ;
	    RECT 143.0000 38.1000 143.3000 38.8000 ;
	    RECT 143.0000 37.8000 151.3000 38.1000 ;
      END
   END OUTPD<3>
   PIN OUTPD<4>
      PORT
         LAYER metal1 ;
	    RECT 142.2000 46.2000 142.6000 49.9000 ;
	    RECT 142.3000 45.1000 142.6000 46.2000 ;
	    RECT 142.2000 41.1000 142.6000 45.1000 ;
         LAYER metal2 ;
	    RECT 142.2000 46.8000 142.6000 47.2000 ;
	    RECT 142.2000 46.2000 142.5000 46.8000 ;
	    RECT 142.2000 45.8000 142.6000 46.2000 ;
         LAYER metal3 ;
	    RECT 142.2000 46.1000 142.6000 46.2000 ;
	    RECT 142.2000 45.8000 151.3000 46.1000 ;
      END
   END OUTPD<4>
   PIN OUTPD<5>
      PORT
         LAYER metal1 ;
	    RECT 144.6000 55.9000 145.0000 59.9000 ;
	    RECT 144.7000 54.8000 145.0000 55.9000 ;
	    RECT 144.6000 51.1000 145.0000 54.8000 ;
         LAYER metal2 ;
	    RECT 144.6000 58.8000 145.0000 59.2000 ;
	    RECT 144.6000 58.2000 144.9000 58.8000 ;
	    RECT 144.6000 57.8000 145.0000 58.2000 ;
         LAYER metal3 ;
	    RECT 144.6000 58.8000 145.0000 59.2000 ;
	    RECT 144.6000 58.1000 144.9000 58.8000 ;
	    RECT 144.6000 57.8000 151.3000 58.1000 ;
      END
   END OUTPD<5>
   PIN OUTPD<6>
      PORT
         LAYER metal1 ;
	    RECT 147.0000 27.1000 147.4000 29.9000 ;
	    RECT 148.6000 27.1000 149.0000 27.2000 ;
	    RECT 147.0000 26.8000 149.0000 27.1000 ;
	    RECT 147.0000 26.2000 147.4000 26.8000 ;
	    RECT 147.1000 25.1000 147.4000 26.2000 ;
	    RECT 147.0000 21.1000 147.4000 25.1000 ;
         LAYER metal2 ;
	    RECT 148.6000 26.8000 149.0000 27.2000 ;
	    RECT 148.6000 26.2000 148.9000 26.8000 ;
	    RECT 148.6000 25.8000 149.0000 26.2000 ;
         LAYER metal3 ;
	    RECT 148.6000 26.1000 149.0000 26.2000 ;
	    RECT 148.6000 25.8000 151.3000 26.1000 ;
      END
   END OUTPD<6>
   PIN OUTPD<7>
      PORT
         LAYER metal1 ;
	    RECT 98.2000 6.2000 98.6000 9.9000 ;
	    RECT 98.3000 5.1000 98.6000 6.2000 ;
	    RECT 98.2000 1.1000 98.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 98.2000 1.8000 98.6000 2.2000 ;
	    RECT 98.2000 -2.2000 98.5000 1.8000 ;
      END
   END OUTPD<7>
   PIN OUTPD<8>
      PORT
         LAYER metal1 ;
	    RECT 0.6000 35.9000 1.0000 39.9000 ;
	    RECT 0.6000 34.8000 0.9000 35.9000 ;
	    RECT 0.6000 31.1000 1.0000 34.8000 ;
         LAYER metal2 ;
	    RECT 0.6000 36.8000 1.0000 37.2000 ;
	    RECT 0.6000 36.2000 0.9000 36.8000 ;
	    RECT 0.6000 35.8000 1.0000 36.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 36.1000 1.0000 36.2000 ;
	    RECT -2.6000 35.8000 1.0000 36.1000 ;
      END
   END OUTPD<8>
   PIN OUTPD<9>
      PORT
         LAYER metal1 ;
	    RECT 101.4000 26.2000 101.8000 29.9000 ;
	    RECT 101.5000 25.1000 101.8000 26.2000 ;
	    RECT 101.4000 21.1000 101.8000 25.1000 ;
         LAYER metal2 ;
	    RECT 101.4000 21.8000 101.8000 22.2000 ;
	    RECT 101.4000 16.2000 101.7000 21.8000 ;
	    RECT 101.4000 15.8000 101.8000 16.2000 ;
	    RECT 102.2000 0.8000 102.6000 1.2000 ;
	    RECT 102.2000 -2.2000 102.5000 0.8000 ;
         LAYER metal3 ;
	    RECT 101.4000 16.1000 101.8000 16.2000 ;
	    RECT 102.2000 16.1000 102.6000 16.2000 ;
	    RECT 101.4000 15.8000 102.6000 16.1000 ;
	    RECT 101.4000 1.1000 101.8000 1.2000 ;
	    RECT 102.2000 1.1000 102.6000 1.2000 ;
	    RECT 101.4000 0.8000 102.6000 1.1000 ;
         LAYER metal4 ;
	    RECT 102.2000 15.8000 102.6000 16.2000 ;
	    RECT 101.4000 1.1000 101.8000 1.2000 ;
	    RECT 102.2000 1.1000 102.5000 15.8000 ;
	    RECT 101.4000 0.8000 102.5000 1.1000 ;
      END
   END OUTPD<9>
   PIN OUTPD<10>
      PORT
         LAYER metal1 ;
	    RECT 0.6000 106.2000 1.0000 109.9000 ;
	    RECT 0.6000 105.1000 0.9000 106.2000 ;
	    RECT 0.6000 101.1000 1.0000 105.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 106.8000 1.0000 107.2000 ;
	    RECT 0.6000 106.2000 0.9000 106.8000 ;
	    RECT 0.6000 105.8000 1.0000 106.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 106.1000 1.0000 106.2000 ;
	    RECT -2.6000 105.8000 1.0000 106.1000 ;
      END
   END OUTPD<10>
   PIN OUTPD<11>
      PORT
         LAYER metal1 ;
	    RECT 137.4000 115.9000 137.8000 119.9000 ;
	    RECT 137.5000 114.8000 137.8000 115.9000 ;
	    RECT 137.4000 111.1000 137.8000 114.8000 ;
         LAYER metal2 ;
	    RECT 137.4000 119.2000 137.7000 123.1000 ;
	    RECT 137.4000 118.8000 137.8000 119.2000 ;
      END
   END OUTPD<11>
   PIN OUTPD<12>
      PORT
         LAYER metal1 ;
	    RECT 0.6000 55.9000 1.0000 59.9000 ;
	    RECT 0.6000 54.8000 0.9000 55.9000 ;
	    RECT 0.6000 51.1000 1.0000 54.8000 ;
         LAYER metal2 ;
	    RECT 0.6000 58.8000 1.0000 59.2000 ;
	    RECT 0.6000 58.2000 0.9000 58.8000 ;
	    RECT 0.6000 57.8000 1.0000 58.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 58.8000 1.0000 59.2000 ;
	    RECT 0.6000 58.1000 0.9000 58.8000 ;
	    RECT -2.6000 57.8000 0.9000 58.1000 ;
      END
   END OUTPD<12>
   PIN OUTPD<13>
      PORT
         LAYER metal1 ;
	    RECT 126.2000 6.2000 126.6000 9.9000 ;
	    RECT 126.3000 5.1000 126.6000 6.2000 ;
	    RECT 126.2000 1.1000 126.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 126.2000 1.8000 126.6000 2.2000 ;
	    RECT 126.2000 -2.2000 126.5000 1.8000 ;
      END
   END OUTPD<13>
   PIN OUTPD<14>
      PORT
         LAYER metal1 ;
	    RECT 86.2000 106.2000 86.6000 109.9000 ;
	    RECT 86.3000 105.1000 86.6000 106.2000 ;
	    RECT 86.2000 101.1000 86.6000 105.1000 ;
         LAYER metal2 ;
	    RECT 86.2000 122.8000 87.3000 123.1000 ;
	    RECT 86.2000 109.2000 86.5000 122.8000 ;
	    RECT 86.2000 108.8000 86.6000 109.2000 ;
      END
   END OUTPD<14>
   PIN OUTPD<15>
      PORT
         LAYER metal1 ;
	    RECT 111.8000 6.2000 112.2000 9.9000 ;
	    RECT 111.9000 5.1000 112.2000 6.2000 ;
	    RECT 111.8000 1.1000 112.2000 5.1000 ;
         LAYER metal2 ;
	    RECT 111.8000 1.8000 112.2000 2.2000 ;
	    RECT 111.8000 -2.2000 112.1000 1.8000 ;
      END
   END OUTPD<15>
   PIN reset
      PORT
         LAYER metal1 ;
	    RECT 0.6000 6.2000 1.0000 9.9000 ;
	    RECT 0.6000 5.1000 0.9000 6.2000 ;
	    RECT 0.6000 1.1000 1.0000 5.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 6.8000 1.0000 7.2000 ;
	    RECT 0.6000 6.2000 0.9000 6.8000 ;
	    RECT 0.6000 5.8000 1.0000 6.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 6.1000 1.0000 6.2000 ;
	    RECT -2.6000 5.8000 1.0000 6.1000 ;
      END
   END reset
   PIN RD
      PORT
         LAYER metal1 ;
	    RECT 79.8000 6.2000 80.2000 9.9000 ;
	    RECT 79.8000 5.1000 80.1000 6.2000 ;
	    RECT 79.8000 1.1000 80.2000 5.1000 ;
         LAYER metal2 ;
	    RECT 79.8000 1.8000 80.2000 2.2000 ;
	    RECT 79.8000 -2.2000 80.1000 1.8000 ;
      END
   END RD
   PIN WD
      PORT
         LAYER metal1 ;
	    RECT 82.2000 6.2000 82.6000 9.9000 ;
	    RECT 82.2000 5.1000 82.5000 6.2000 ;
	    RECT 82.2000 1.1000 82.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 82.2000 1.8000 82.6000 2.2000 ;
	    RECT 82.2000 -2.2000 82.5000 1.8000 ;
      END
   END WD
   PIN WDATA<0>
      PORT
         LAYER metal1 ;
	    RECT 103.8000 26.2000 104.2000 29.9000 ;
	    RECT 103.9000 25.1000 104.2000 26.2000 ;
	    RECT 103.8000 21.1000 104.2000 25.1000 ;
         LAYER metal2 ;
	    RECT 103.8000 21.8000 104.2000 22.2000 ;
	    RECT 103.8000 14.1000 104.1000 21.8000 ;
	    RECT 104.6000 14.1000 105.0000 14.2000 ;
	    RECT 103.8000 13.8000 105.0000 14.1000 ;
	    RECT 103.8000 0.8000 104.2000 1.2000 ;
	    RECT 103.8000 -2.2000 104.1000 0.8000 ;
         LAYER metal3 ;
	    RECT 103.8000 14.1000 104.2000 14.2000 ;
	    RECT 104.6000 14.1000 105.0000 14.2000 ;
	    RECT 103.8000 13.8000 105.0000 14.1000 ;
	    RECT 103.8000 1.8000 104.2000 2.2000 ;
	    RECT 103.8000 1.2000 104.1000 1.8000 ;
	    RECT 103.8000 0.8000 104.2000 1.2000 ;
         LAYER metal4 ;
	    RECT 103.8000 13.8000 104.2000 14.2000 ;
	    RECT 103.8000 2.2000 104.1000 13.8000 ;
	    RECT 103.8000 1.8000 104.2000 2.2000 ;
      END
   END WDATA<0>
   PIN WDATA<1>
      PORT
         LAYER metal1 ;
	    RECT 94.2000 115.9000 94.6000 119.9000 ;
	    RECT 94.3000 114.8000 94.6000 115.9000 ;
	    RECT 94.2000 111.1000 94.6000 114.8000 ;
         LAYER metal2 ;
	    RECT 94.2000 122.8000 95.3000 123.1000 ;
	    RECT 94.2000 119.2000 94.5000 122.8000 ;
	    RECT 94.2000 118.8000 94.6000 119.2000 ;
      END
   END WDATA<1>
   PIN WDATA<2>
      PORT
         LAYER metal1 ;
	    RECT 99.8000 95.9000 100.2000 99.9000 ;
	    RECT 99.8000 94.8000 100.1000 95.9000 ;
	    RECT 99.8000 91.1000 100.2000 94.8000 ;
         LAYER metal2 ;
	    RECT 99.8000 121.2000 100.1000 123.1000 ;
	    RECT 99.8000 120.8000 100.2000 121.2000 ;
	    RECT 99.8000 100.8000 100.2000 101.2000 ;
	    RECT 99.8000 99.2000 100.1000 100.8000 ;
	    RECT 99.8000 98.8000 100.2000 99.2000 ;
         LAYER metal3 ;
	    RECT 99.8000 120.8000 100.2000 121.2000 ;
	    RECT 99.8000 120.2000 100.1000 120.8000 ;
	    RECT 99.8000 119.8000 100.2000 120.2000 ;
	    RECT 99.8000 101.8000 100.2000 102.2000 ;
	    RECT 99.8000 101.2000 100.1000 101.8000 ;
	    RECT 99.8000 100.8000 100.2000 101.2000 ;
         LAYER metal4 ;
	    RECT 99.8000 119.8000 100.2000 120.2000 ;
	    RECT 99.8000 102.2000 100.1000 119.8000 ;
	    RECT 99.8000 101.8000 100.2000 102.2000 ;
      END
   END WDATA<2>
   PIN WDATA<3>
      PORT
         LAYER metal1 ;
	    RECT 139.8000 55.9000 140.2000 59.9000 ;
	    RECT 139.9000 54.8000 140.2000 55.9000 ;
	    RECT 139.8000 51.1000 140.2000 54.8000 ;
         LAYER metal2 ;
	    RECT 139.8000 57.8000 140.2000 58.2000 ;
	    RECT 139.8000 57.2000 140.1000 57.8000 ;
	    RECT 139.8000 56.8000 140.2000 57.2000 ;
         LAYER metal3 ;
	    RECT 139.8000 57.8000 140.2000 58.2000 ;
	    RECT 139.8000 57.1000 140.1000 57.8000 ;
	    RECT 139.8000 56.8000 151.3000 57.1000 ;
	    RECT 151.0000 55.8000 151.3000 56.8000 ;
      END
   END WDATA<3>
   PIN WDATA<4>
      PORT
         LAYER metal1 ;
	    RECT 145.4000 79.1000 145.8000 79.9000 ;
	    RECT 148.6000 79.1000 149.0000 79.2000 ;
	    RECT 145.4000 78.8000 149.0000 79.1000 ;
	    RECT 145.4000 75.9000 145.8000 78.8000 ;
	    RECT 145.5000 74.8000 145.8000 75.9000 ;
	    RECT 145.4000 71.1000 145.8000 74.8000 ;
         LAYER metal2 ;
	    RECT 148.6000 79.8000 149.0000 80.2000 ;
	    RECT 148.6000 79.2000 148.9000 79.8000 ;
	    RECT 148.6000 78.8000 149.0000 79.2000 ;
         LAYER metal3 ;
	    RECT 148.6000 80.1000 149.0000 80.2000 ;
	    RECT 148.6000 79.8000 151.3000 80.1000 ;
      END
   END WDATA<4>
   PIN WDATA<5>
      PORT
         LAYER metal1 ;
	    RECT 106.2000 115.9000 106.6000 119.9000 ;
	    RECT 106.3000 114.8000 106.6000 115.9000 ;
	    RECT 106.2000 111.1000 106.6000 114.8000 ;
         LAYER metal2 ;
	    RECT 107.8000 121.2000 108.1000 123.1000 ;
	    RECT 106.2000 120.8000 106.6000 121.2000 ;
	    RECT 107.8000 120.8000 108.2000 121.2000 ;
	    RECT 106.2000 119.2000 106.5000 120.8000 ;
	    RECT 106.2000 118.8000 106.6000 119.2000 ;
         LAYER metal3 ;
	    RECT 106.2000 121.1000 106.6000 121.2000 ;
	    RECT 107.8000 121.1000 108.2000 121.2000 ;
	    RECT 106.2000 120.8000 108.2000 121.1000 ;
      END
   END WDATA<5>
   PIN WDATA<6>
      PORT
         LAYER metal1 ;
	    RECT 142.2000 95.9000 142.6000 99.9000 ;
	    RECT 142.3000 94.8000 142.6000 95.9000 ;
	    RECT 142.2000 91.1000 142.6000 94.8000 ;
         LAYER metal2 ;
	    RECT 142.2000 98.8000 142.6000 99.2000 ;
	    RECT 142.2000 98.2000 142.5000 98.8000 ;
	    RECT 142.2000 97.8000 142.6000 98.2000 ;
         LAYER metal3 ;
	    RECT 142.2000 98.8000 142.6000 99.2000 ;
	    RECT 142.2000 98.1000 142.5000 98.8000 ;
	    RECT 142.2000 97.8000 151.3000 98.1000 ;
      END
   END WDATA<6>
   PIN WDATA<7>
      PORT
         LAYER metal1 ;
	    RECT 147.0000 87.1000 147.4000 89.9000 ;
	    RECT 148.6000 87.1000 149.0000 87.2000 ;
	    RECT 147.0000 86.8000 149.0000 87.1000 ;
	    RECT 147.0000 86.2000 147.4000 86.8000 ;
	    RECT 147.1000 85.1000 147.4000 86.2000 ;
	    RECT 147.0000 81.1000 147.4000 85.1000 ;
         LAYER metal2 ;
	    RECT 148.6000 86.8000 149.0000 87.2000 ;
	    RECT 148.6000 86.2000 148.9000 86.8000 ;
	    RECT 148.6000 85.8000 149.0000 86.2000 ;
         LAYER metal3 ;
	    RECT 148.6000 86.1000 149.0000 86.2000 ;
	    RECT 148.6000 85.8000 151.3000 86.1000 ;
      END
   END WDATA<7>
   PIN DP<0>
      PORT
         LAYER metal1 ;
	    RECT 0.6000 75.9000 1.0000 79.9000 ;
	    RECT 0.6000 74.8000 0.9000 75.9000 ;
	    RECT 0.6000 71.1000 1.0000 74.8000 ;
         LAYER metal2 ;
	    RECT 0.6000 76.8000 1.0000 77.2000 ;
	    RECT 0.6000 76.2000 0.9000 76.8000 ;
	    RECT 0.6000 75.8000 1.0000 76.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 76.1000 1.0000 76.2000 ;
	    RECT -2.6000 75.8000 1.0000 76.1000 ;
      END
   END DP<0>
   PIN DP<1>
      PORT
         LAYER metal1 ;
	    RECT 0.6000 95.9000 1.0000 99.9000 ;
	    RECT 0.6000 94.8000 0.9000 95.9000 ;
	    RECT 0.6000 91.1000 1.0000 94.8000 ;
         LAYER metal2 ;
	    RECT 0.6000 98.8000 1.0000 99.2000 ;
	    RECT 0.6000 98.2000 0.9000 98.8000 ;
	    RECT 0.6000 97.8000 1.0000 98.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 98.8000 1.0000 99.2000 ;
	    RECT 0.6000 98.1000 0.9000 98.8000 ;
	    RECT -2.6000 97.8000 0.9000 98.1000 ;
      END
   END DP<1>
   PIN DP<2>
      PORT
         LAYER metal1 ;
	    RECT 3.0000 95.9000 3.4000 99.9000 ;
	    RECT 3.0000 94.8000 3.3000 95.9000 ;
	    RECT 3.0000 91.1000 3.4000 94.8000 ;
         LAYER metal2 ;
	    RECT 3.0000 96.8000 3.4000 97.2000 ;
	    RECT 3.0000 96.2000 3.3000 96.8000 ;
	    RECT 3.0000 95.8000 3.4000 96.2000 ;
         LAYER metal3 ;
	    RECT 3.0000 96.1000 3.4000 96.2000 ;
	    RECT -2.6000 95.8000 3.4000 96.1000 ;
      END
   END DP<2>
   PIN DP<3>
      PORT
         LAYER metal1 ;
	    RECT 0.6000 66.2000 1.0000 69.9000 ;
	    RECT 0.6000 65.1000 0.9000 66.2000 ;
	    RECT 0.6000 61.1000 1.0000 65.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 66.8000 1.0000 67.2000 ;
	    RECT 0.6000 66.2000 0.9000 66.8000 ;
	    RECT 0.6000 65.8000 1.0000 66.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 66.1000 1.0000 66.2000 ;
	    RECT -2.6000 65.8000 1.0000 66.1000 ;
      END
   END DP<3>
   PIN DP<4>
      PORT
         LAYER metal1 ;
	    RECT 61.4000 46.2000 61.8000 49.9000 ;
	    RECT 61.5000 45.1000 61.8000 46.2000 ;
	    RECT 61.4000 41.1000 61.8000 45.1000 ;
         LAYER metal2 ;
	    RECT 61.4000 41.8000 61.8000 42.2000 ;
	    RECT 61.4000 37.2000 61.7000 41.8000 ;
	    RECT 61.4000 36.8000 61.8000 37.2000 ;
	    RECT 63.0000 0.8000 63.4000 1.2000 ;
	    RECT 63.0000 -2.2000 63.3000 0.8000 ;
         LAYER metal3 ;
	    RECT 61.4000 37.1000 61.8000 37.2000 ;
	    RECT 63.0000 37.1000 63.4000 37.2000 ;
	    RECT 61.4000 36.8000 63.4000 37.1000 ;
	    RECT 62.2000 1.1000 62.6000 1.2000 ;
	    RECT 63.0000 1.1000 63.4000 1.2000 ;
	    RECT 62.2000 0.8000 63.4000 1.1000 ;
         LAYER metal4 ;
	    RECT 63.0000 36.8000 63.4000 37.2000 ;
	    RECT 62.2000 1.1000 62.6000 1.2000 ;
	    RECT 63.0000 1.1000 63.3000 36.8000 ;
	    RECT 62.2000 0.8000 63.3000 1.1000 ;
      END
   END DP<4>
   PIN DP<5>
      PORT
         LAYER metal1 ;
	    RECT 59.0000 46.2000 59.4000 49.9000 ;
	    RECT 59.1000 45.1000 59.4000 46.2000 ;
	    RECT 59.0000 41.1000 59.4000 45.1000 ;
         LAYER metal2 ;
	    RECT 59.0000 41.8000 59.4000 42.2000 ;
	    RECT 59.0000 27.2000 59.3000 41.8000 ;
	    RECT 59.0000 26.8000 59.4000 27.2000 ;
	    RECT 59.0000 0.8000 59.4000 1.2000 ;
	    RECT 59.0000 -2.2000 59.3000 0.8000 ;
         LAYER metal3 ;
	    RECT 58.2000 27.1000 58.6000 27.2000 ;
	    RECT 59.0000 27.1000 59.4000 27.2000 ;
	    RECT 58.2000 26.8000 59.4000 27.1000 ;
	    RECT 59.0000 1.8000 59.4000 2.2000 ;
	    RECT 59.0000 1.2000 59.3000 1.8000 ;
	    RECT 59.0000 0.8000 59.4000 1.2000 ;
         LAYER metal4 ;
	    RECT 58.2000 27.1000 58.6000 27.2000 ;
	    RECT 58.2000 26.8000 59.3000 27.1000 ;
	    RECT 59.0000 2.2000 59.3000 26.8000 ;
	    RECT 59.0000 1.8000 59.4000 2.2000 ;
      END
   END DP<5>
   PIN DP<6>
      PORT
         LAYER metal1 ;
	    RECT 84.6000 115.9000 85.0000 119.9000 ;
	    RECT 84.7000 114.8000 85.0000 115.9000 ;
	    RECT 84.6000 111.1000 85.0000 114.8000 ;
         LAYER metal2 ;
	    RECT 84.6000 119.2000 84.9000 123.1000 ;
	    RECT 84.6000 118.8000 85.0000 119.2000 ;
      END
   END DP<6>
   PIN DP<7>
      PORT
         LAYER metal1 ;
	    RECT 61.4000 95.9000 61.8000 99.9000 ;
	    RECT 61.5000 94.8000 61.8000 95.9000 ;
	    RECT 61.4000 91.1000 61.8000 94.8000 ;
         LAYER metal2 ;
	    RECT 61.4000 121.2000 61.7000 123.1000 ;
	    RECT 61.4000 120.8000 61.8000 121.2000 ;
	    RECT 61.4000 103.8000 61.8000 104.2000 ;
	    RECT 61.4000 99.2000 61.7000 103.8000 ;
	    RECT 61.4000 98.8000 61.8000 99.2000 ;
         LAYER metal3 ;
	    RECT 61.4000 120.8000 61.8000 121.2000 ;
	    RECT 61.4000 120.2000 61.7000 120.8000 ;
	    RECT 61.4000 119.8000 61.8000 120.2000 ;
	    RECT 61.4000 104.8000 61.8000 105.2000 ;
	    RECT 61.4000 104.2000 61.7000 104.8000 ;
	    RECT 61.4000 103.8000 61.8000 104.2000 ;
         LAYER metal4 ;
	    RECT 61.4000 119.8000 61.8000 120.2000 ;
	    RECT 61.4000 105.2000 61.7000 119.8000 ;
	    RECT 61.4000 104.8000 61.8000 105.2000 ;
      END
   END DP<7>
   PIN DP<8>
      PORT
         LAYER metal1 ;
	    RECT 0.6000 86.2000 1.0000 89.9000 ;
	    RECT 0.6000 85.1000 0.9000 86.2000 ;
	    RECT 0.6000 81.1000 1.0000 85.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 86.8000 1.0000 87.2000 ;
	    RECT 0.6000 86.2000 0.9000 86.8000 ;
	    RECT 0.6000 85.8000 1.0000 86.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 86.1000 1.0000 86.2000 ;
	    RECT -2.6000 85.8000 1.0000 86.1000 ;
      END
   END DP<8>
   PIN DP<9>
      PORT
         LAYER metal1 ;
	    RECT 47.8000 119.1000 48.2000 119.9000 ;
	    RECT 49.4000 119.1000 49.8000 119.2000 ;
	    RECT 47.8000 118.8000 49.8000 119.1000 ;
	    RECT 47.8000 115.9000 48.2000 118.8000 ;
	    RECT 47.9000 114.8000 48.2000 115.9000 ;
	    RECT 47.8000 111.1000 48.2000 114.8000 ;
         LAYER metal2 ;
	    RECT 47.8000 122.8000 49.7000 123.1000 ;
	    RECT 49.4000 119.2000 49.7000 122.8000 ;
	    RECT 49.4000 118.8000 49.8000 119.2000 ;
      END
   END DP<9>
   PIN DP<10>
      PORT
         LAYER metal1 ;
	    RECT 16.6000 106.2000 17.0000 109.9000 ;
	    RECT 16.6000 105.1000 16.9000 106.2000 ;
	    RECT 16.6000 101.1000 17.0000 105.1000 ;
         LAYER metal2 ;
	    RECT 16.6000 121.2000 16.9000 123.1000 ;
	    RECT 16.6000 120.8000 17.0000 121.2000 ;
	    RECT 16.6000 110.8000 17.0000 111.2000 ;
	    RECT 16.6000 109.2000 16.9000 110.8000 ;
	    RECT 16.6000 108.8000 17.0000 109.2000 ;
         LAYER metal3 ;
	    RECT 16.6000 120.8000 17.0000 121.2000 ;
	    RECT 16.6000 120.2000 16.9000 120.8000 ;
	    RECT 16.6000 119.8000 17.0000 120.2000 ;
	    RECT 16.6000 111.8000 17.0000 112.2000 ;
	    RECT 16.6000 111.2000 16.9000 111.8000 ;
	    RECT 16.6000 110.8000 17.0000 111.2000 ;
         LAYER metal4 ;
	    RECT 16.6000 119.8000 17.0000 120.2000 ;
	    RECT 16.6000 112.2000 16.9000 119.8000 ;
	    RECT 16.6000 111.8000 17.0000 112.2000 ;
      END
   END DP<10>
   PIN DP<11>
      PORT
         LAYER metal1 ;
	    RECT 10.2000 115.9000 10.6000 119.9000 ;
	    RECT 10.2000 114.8000 10.5000 115.9000 ;
	    RECT 10.2000 111.1000 10.6000 114.8000 ;
         LAYER metal2 ;
	    RECT 10.2000 119.2000 10.5000 123.1000 ;
	    RECT 10.2000 118.8000 10.6000 119.2000 ;
      END
   END DP<11>
   PIN DP<12>
      PORT
         LAYER metal1 ;
	    RECT 82.2000 115.9000 82.6000 119.9000 ;
	    RECT 82.3000 114.8000 82.6000 115.9000 ;
	    RECT 82.2000 111.1000 82.6000 114.8000 ;
         LAYER metal2 ;
	    RECT 82.2000 119.2000 82.5000 123.1000 ;
	    RECT 82.2000 118.8000 82.6000 119.2000 ;
      END
   END DP<12>
   PIN DP<13>
      PORT
         LAYER metal1 ;
	    RECT 70.2000 115.9000 70.6000 119.9000 ;
	    RECT 70.3000 114.8000 70.6000 115.9000 ;
	    RECT 70.2000 111.1000 70.6000 114.8000 ;
         LAYER metal2 ;
	    RECT 70.2000 119.2000 70.5000 123.1000 ;
	    RECT 70.2000 118.8000 70.6000 119.2000 ;
      END
   END DP<13>
   PIN DP<14>
      PORT
         LAYER metal1 ;
	    RECT 21.4000 115.9000 21.8000 119.9000 ;
	    RECT 21.5000 114.8000 21.8000 115.9000 ;
	    RECT 21.4000 111.1000 21.8000 114.8000 ;
         LAYER metal2 ;
	    RECT 21.4000 119.2000 21.7000 123.1000 ;
	    RECT 21.4000 118.8000 21.8000 119.2000 ;
      END
   END DP<14>
   PIN PCDELTA<0>
      PORT
         LAYER metal1 ;
	    RECT 66.2000 6.2000 66.6000 9.9000 ;
	    RECT 66.3000 5.1000 66.6000 6.2000 ;
	    RECT 66.2000 1.1000 66.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 66.2000 1.8000 66.6000 2.2000 ;
	    RECT 66.2000 -2.2000 66.5000 1.8000 ;
      END
   END PCDELTA<0>
   PIN PCDELTA<1>
      PORT
         LAYER metal1 ;
	    RECT 3.0000 55.9000 3.4000 59.9000 ;
	    RECT 3.0000 54.8000 3.3000 55.9000 ;
	    RECT 3.0000 51.1000 3.4000 54.8000 ;
         LAYER metal2 ;
	    RECT 3.0000 56.8000 3.4000 57.2000 ;
	    RECT 3.0000 56.2000 3.3000 56.8000 ;
	    RECT 3.0000 55.8000 3.4000 56.2000 ;
         LAYER metal3 ;
	    RECT 3.0000 56.1000 3.4000 56.2000 ;
	    RECT -2.6000 55.8000 3.4000 56.1000 ;
      END
   END PCDELTA<1>
   PIN PCDELTA<2>
      PORT
         LAYER metal1 ;
	    RECT 144.6000 115.9000 145.0000 119.9000 ;
	    RECT 144.7000 114.8000 145.0000 115.9000 ;
	    RECT 144.6000 111.1000 145.0000 114.8000 ;
         LAYER metal2 ;
	    RECT 144.6000 119.2000 144.9000 123.1000 ;
	    RECT 144.6000 118.8000 145.0000 119.2000 ;
      END
   END PCDELTA<2>
   PIN PCDELTA<3>
      PORT
         LAYER metal1 ;
	    RECT 89.4000 115.9000 89.8000 119.9000 ;
	    RECT 89.5000 114.8000 89.8000 115.9000 ;
	    RECT 89.4000 111.1000 89.8000 114.8000 ;
         LAYER metal2 ;
	    RECT 91.0000 121.2000 91.3000 123.1000 ;
	    RECT 89.4000 120.8000 89.8000 121.2000 ;
	    RECT 91.0000 120.8000 91.4000 121.2000 ;
	    RECT 89.4000 119.2000 89.7000 120.8000 ;
	    RECT 89.4000 118.8000 89.8000 119.2000 ;
         LAYER metal3 ;
	    RECT 89.4000 121.1000 89.8000 121.2000 ;
	    RECT 91.0000 121.1000 91.4000 121.2000 ;
	    RECT 89.4000 120.8000 91.4000 121.1000 ;
      END
   END PCDELTA<3>
   PIN PCDELTA<4>
      PORT
         LAYER metal1 ;
	    RECT 114.2000 6.2000 114.6000 9.9000 ;
	    RECT 114.3000 5.1000 114.6000 6.2000 ;
	    RECT 114.2000 1.1000 114.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 114.2000 1.8000 114.6000 2.2000 ;
	    RECT 114.2000 -2.2000 114.5000 1.8000 ;
      END
   END PCDELTA<4>
   PIN PCDELTA<5>
      PORT
         LAYER metal1 ;
	    RECT 91.8000 115.9000 92.2000 119.9000 ;
	    RECT 91.9000 114.8000 92.2000 115.9000 ;
	    RECT 91.8000 111.1000 92.2000 114.8000 ;
         LAYER metal2 ;
	    RECT 93.4000 121.2000 93.7000 123.1000 ;
	    RECT 91.8000 120.8000 92.2000 121.2000 ;
	    RECT 93.4000 120.8000 93.8000 121.2000 ;
	    RECT 91.8000 119.2000 92.1000 120.8000 ;
	    RECT 91.8000 118.8000 92.2000 119.2000 ;
         LAYER metal3 ;
	    RECT 91.8000 121.1000 92.2000 121.2000 ;
	    RECT 93.4000 121.1000 93.8000 121.2000 ;
	    RECT 91.8000 120.8000 93.8000 121.1000 ;
      END
   END PCDELTA<5>
   PIN PCDELTA<6>
      PORT
         LAYER metal1 ;
	    RECT 139.0000 6.2000 139.4000 9.9000 ;
	    RECT 139.1000 5.1000 139.4000 6.2000 ;
	    RECT 139.0000 1.1000 139.4000 5.1000 ;
         LAYER metal2 ;
	    RECT 139.0000 1.8000 139.4000 2.2000 ;
	    RECT 139.0000 -2.2000 139.3000 1.8000 ;
      END
   END PCDELTA<6>
   PIN PCDELTA<7>
      PORT
         LAYER metal1 ;
	    RECT 145.4000 37.1000 145.8000 39.9000 ;
	    RECT 148.6000 37.1000 149.0000 37.2000 ;
	    RECT 145.4000 36.8000 149.0000 37.1000 ;
	    RECT 145.4000 35.9000 145.8000 36.8000 ;
	    RECT 145.5000 34.8000 145.8000 35.9000 ;
	    RECT 145.4000 31.1000 145.8000 34.8000 ;
         LAYER metal2 ;
	    RECT 148.6000 36.8000 149.0000 37.2000 ;
	    RECT 148.6000 36.2000 148.9000 36.8000 ;
	    RECT 148.6000 35.8000 149.0000 36.2000 ;
         LAYER metal3 ;
	    RECT 148.6000 36.1000 149.0000 36.2000 ;
	    RECT 148.6000 35.8000 151.3000 36.1000 ;
      END
   END PCDELTA<7>
   PIN PCDELTA<8>
      PORT
         LAYER metal1 ;
	    RECT 143.8000 6.2000 144.2000 9.9000 ;
	    RECT 143.9000 5.1000 144.2000 6.2000 ;
	    RECT 143.8000 1.1000 144.2000 5.1000 ;
         LAYER metal2 ;
	    RECT 143.8000 1.8000 144.2000 2.2000 ;
	    RECT 143.8000 -2.2000 144.1000 1.8000 ;
      END
   END PCDELTA<8>
   PIN PCDELTA<9>
      PORT
         LAYER metal1 ;
	    RECT 141.4000 6.2000 141.8000 9.9000 ;
	    RECT 141.5000 5.1000 141.8000 6.2000 ;
	    RECT 141.4000 1.1000 141.8000 5.1000 ;
         LAYER metal2 ;
	    RECT 141.4000 1.8000 141.8000 2.2000 ;
	    RECT 141.4000 -2.2000 141.7000 1.8000 ;
      END
   END PCDELTA<9>
   PIN PCDELTA<10>
      PORT
         LAYER metal1 ;
	    RECT 146.2000 99.1000 146.6000 99.9000 ;
	    RECT 148.6000 99.1000 149.0000 99.2000 ;
	    RECT 146.2000 98.8000 149.0000 99.1000 ;
	    RECT 146.2000 95.9000 146.6000 98.8000 ;
	    RECT 146.3000 94.8000 146.6000 95.9000 ;
	    RECT 146.2000 91.1000 146.6000 94.8000 ;
         LAYER metal2 ;
	    RECT 148.6000 99.8000 149.0000 100.2000 ;
	    RECT 148.6000 99.2000 148.9000 99.8000 ;
	    RECT 148.6000 98.8000 149.0000 99.2000 ;
         LAYER metal3 ;
	    RECT 148.6000 100.1000 149.0000 100.2000 ;
	    RECT 148.6000 99.8000 151.3000 100.1000 ;
      END
   END PCDELTA<10>
   PIN PCDELTA<11>
      PORT
         LAYER metal1 ;
	    RECT 142.2000 115.9000 142.6000 119.9000 ;
	    RECT 142.3000 114.8000 142.6000 115.9000 ;
	    RECT 142.2000 111.1000 142.6000 114.8000 ;
         LAYER metal2 ;
	    RECT 142.2000 119.2000 142.5000 123.1000 ;
	    RECT 142.2000 118.8000 142.6000 119.2000 ;
      END
   END PCDELTA<11>
   PIN PCDELTA<12>
      PORT
         LAYER metal1 ;
	    RECT 121.4000 6.2000 121.8000 9.9000 ;
	    RECT 121.5000 5.1000 121.8000 6.2000 ;
	    RECT 121.4000 1.1000 121.8000 5.1000 ;
         LAYER metal2 ;
	    RECT 121.4000 1.8000 121.8000 2.2000 ;
	    RECT 121.4000 -2.2000 121.7000 1.8000 ;
      END
   END PCDELTA<12>
   PIN PCDELTA<13>
      PORT
         LAYER metal1 ;
	    RECT 147.0000 69.1000 147.4000 69.9000 ;
	    RECT 148.6000 69.1000 149.0000 69.2000 ;
	    RECT 147.0000 68.8000 149.0000 69.1000 ;
	    RECT 147.0000 66.2000 147.4000 68.8000 ;
	    RECT 147.1000 65.1000 147.4000 66.2000 ;
	    RECT 147.0000 61.1000 147.4000 65.1000 ;
         LAYER metal2 ;
	    RECT 148.6000 69.8000 149.0000 70.2000 ;
	    RECT 148.6000 69.2000 148.9000 69.8000 ;
	    RECT 148.6000 68.8000 149.0000 69.2000 ;
         LAYER metal3 ;
	    RECT 148.6000 70.1000 149.0000 70.2000 ;
	    RECT 148.6000 69.8000 151.3000 70.1000 ;
      END
   END PCDELTA<13>
   PIN PCDELTA<14>
      PORT
         LAYER metal1 ;
	    RECT 147.0000 117.1000 147.4000 119.9000 ;
	    RECT 148.6000 117.1000 149.0000 117.2000 ;
	    RECT 147.0000 116.8000 149.0000 117.1000 ;
	    RECT 147.0000 115.9000 147.4000 116.8000 ;
	    RECT 147.1000 114.8000 147.4000 115.9000 ;
	    RECT 147.0000 111.1000 147.4000 114.8000 ;
         LAYER metal2 ;
	    RECT 148.6000 116.8000 149.0000 117.2000 ;
	    RECT 148.6000 116.2000 148.9000 116.8000 ;
	    RECT 148.6000 115.8000 149.0000 116.2000 ;
         LAYER metal3 ;
	    RECT 148.6000 116.1000 149.0000 116.2000 ;
	    RECT 148.6000 115.8000 151.3000 116.1000 ;
      END
   END PCDELTA<14>
   PIN PCDELTA<15>
      PORT
         LAYER metal1 ;
	    RECT 87.0000 115.9000 87.4000 119.9000 ;
	    RECT 87.1000 114.8000 87.4000 115.9000 ;
	    RECT 87.0000 111.1000 87.4000 114.8000 ;
         LAYER metal2 ;
	    RECT 88.6000 122.8000 89.7000 123.1000 ;
	    RECT 88.6000 121.2000 88.9000 122.8000 ;
	    RECT 87.0000 120.8000 87.4000 121.2000 ;
	    RECT 88.6000 120.8000 89.0000 121.2000 ;
	    RECT 87.0000 119.2000 87.3000 120.8000 ;
	    RECT 87.0000 118.8000 87.4000 119.2000 ;
         LAYER metal3 ;
	    RECT 87.0000 121.1000 87.4000 121.2000 ;
	    RECT 88.6000 121.1000 89.0000 121.2000 ;
	    RECT 87.0000 120.8000 89.0000 121.1000 ;
      END
   END PCDELTA<15>
   OBS
         LAYER metal1 ;
	    RECT 0.6000 115.6000 1.0000 119.9000 ;
	    RECT 2.7000 117.9000 3.3000 119.9000 ;
	    RECT 5.0000 117.9000 5.4000 119.9000 ;
	    RECT 7.2000 118.2000 7.6000 119.9000 ;
	    RECT 7.2000 117.9000 8.2000 118.2000 ;
	    RECT 3.0000 117.5000 3.4000 117.9000 ;
	    RECT 5.1000 117.6000 5.4000 117.9000 ;
	    RECT 4.7000 117.3000 6.5000 117.6000 ;
	    RECT 7.8000 117.5000 8.2000 117.9000 ;
	    RECT 4.7000 117.2000 5.1000 117.3000 ;
	    RECT 6.1000 117.2000 6.5000 117.3000 ;
	    RECT 2.6000 116.6000 3.3000 117.0000 ;
	    RECT 3.0000 116.1000 3.3000 116.6000 ;
	    RECT 4.1000 116.5000 5.2000 116.8000 ;
	    RECT 4.1000 116.4000 4.5000 116.5000 ;
	    RECT 3.0000 115.8000 4.2000 116.1000 ;
	    RECT 0.6000 115.3000 2.7000 115.6000 ;
	    RECT 0.6000 113.6000 1.0000 115.3000 ;
	    RECT 2.3000 115.2000 2.7000 115.3000 ;
	    RECT 1.5000 114.9000 1.9000 115.0000 ;
	    RECT 1.5000 114.6000 3.4000 114.9000 ;
	    RECT 3.0000 114.5000 3.4000 114.6000 ;
	    RECT 3.9000 114.2000 4.2000 115.8000 ;
	    RECT 4.9000 115.9000 5.2000 116.5000 ;
	    RECT 5.5000 116.5000 5.9000 116.6000 ;
	    RECT 7.8000 116.5000 8.2000 116.6000 ;
	    RECT 5.5000 116.2000 8.2000 116.5000 ;
	    RECT 4.9000 115.7000 7.3000 115.9000 ;
	    RECT 9.4000 115.7000 9.8000 119.9000 ;
	    RECT 11.8000 116.2000 12.2000 119.9000 ;
	    RECT 4.9000 115.6000 9.8000 115.7000 ;
	    RECT 11.1000 115.9000 12.2000 116.2000 ;
	    RECT 12.6000 116.2000 13.0000 119.9000 ;
	    RECT 13.4000 116.2000 13.8000 116.3000 ;
	    RECT 14.8000 116.2000 15.6000 119.9000 ;
	    RECT 12.6000 115.9000 13.8000 116.2000 ;
	    RECT 14.6000 115.9000 15.6000 116.2000 ;
	    RECT 16.7000 116.2000 17.1000 116.3000 ;
	    RECT 17.4000 116.2000 17.8000 119.9000 ;
	    RECT 16.7000 115.9000 17.8000 116.2000 ;
	    RECT 11.1000 115.6000 11.4000 115.9000 ;
	    RECT 6.9000 115.5000 9.8000 115.6000 ;
	    RECT 7.0000 115.4000 9.8000 115.5000 ;
	    RECT 10.8000 115.2000 11.4000 115.6000 ;
	    RECT 14.6000 115.2000 14.9000 115.9000 ;
	    RECT 16.7000 115.6000 17.0000 115.9000 ;
	    RECT 15.3000 115.3000 17.0000 115.6000 ;
	    RECT 15.3000 115.2000 15.7000 115.3000 ;
	    RECT 6.2000 115.1000 6.6000 115.2000 ;
	    RECT 6.2000 114.8000 8.7000 115.1000 ;
	    RECT 7.0000 114.7000 7.4000 114.8000 ;
	    RECT 8.3000 114.7000 8.7000 114.8000 ;
	    RECT 7.5000 114.2000 7.9000 114.3000 ;
	    RECT 3.9000 113.9000 9.4000 114.2000 ;
	    RECT 4.1000 113.8000 4.5000 113.9000 ;
	    RECT 0.6000 113.3000 2.5000 113.6000 ;
	    RECT 0.6000 111.1000 1.0000 113.3000 ;
	    RECT 2.1000 113.2000 2.5000 113.3000 ;
	    RECT 7.0000 113.2000 7.3000 113.9000 ;
	    RECT 8.6000 113.8000 9.4000 113.9000 ;
	    RECT 11.1000 113.7000 11.4000 115.2000 ;
	    RECT 11.8000 115.1000 12.2000 115.2000 ;
	    RECT 11.8000 114.8000 12.9000 115.1000 ;
	    RECT 14.2000 114.9000 14.9000 115.2000 ;
	    RECT 16.4000 114.9000 16.8000 115.0000 ;
	    RECT 14.2000 114.8000 15.1000 114.9000 ;
	    RECT 11.8000 114.4000 12.2000 114.8000 ;
	    RECT 12.6000 114.2000 12.9000 114.8000 ;
	    RECT 14.6000 114.6000 15.1000 114.8000 ;
	    RECT 12.6000 113.8000 13.4000 114.2000 ;
	    RECT 14.0000 113.8000 14.4000 114.2000 ;
	    RECT 6.1000 112.7000 6.5000 112.8000 ;
	    RECT 3.0000 112.1000 3.4000 112.5000 ;
	    RECT 5.1000 112.4000 6.5000 112.7000 ;
	    RECT 7.0000 112.4000 7.4000 113.2000 ;
	    RECT 5.1000 112.1000 5.4000 112.4000 ;
	    RECT 7.8000 112.1000 8.2000 112.5000 ;
	    RECT 2.7000 111.8000 3.4000 112.1000 ;
	    RECT 2.7000 111.1000 3.3000 111.8000 ;
	    RECT 5.0000 111.1000 5.4000 112.1000 ;
	    RECT 7.2000 111.8000 8.2000 112.1000 ;
	    RECT 7.2000 111.1000 7.6000 111.8000 ;
	    RECT 9.4000 111.1000 9.8000 113.5000 ;
	    RECT 11.1000 113.4000 12.2000 113.7000 ;
	    RECT 14.1000 113.6000 14.4000 113.8000 ;
	    RECT 13.4000 113.4000 13.8000 113.5000 ;
	    RECT 11.8000 111.1000 12.2000 113.4000 ;
	    RECT 12.6000 113.1000 13.8000 113.4000 ;
	    RECT 14.1000 113.2000 14.5000 113.6000 ;
	    RECT 12.6000 111.1000 13.0000 113.1000 ;
	    RECT 14.8000 112.9000 15.1000 114.6000 ;
	    RECT 15.5000 114.6000 16.8000 114.9000 ;
	    RECT 15.5000 114.3000 15.8000 114.6000 ;
	    RECT 15.4000 113.9000 15.8000 114.3000 ;
	    RECT 17.0000 114.1000 17.8000 114.2000 ;
	    RECT 16.1000 113.8000 17.8000 114.1000 ;
	    RECT 16.1000 113.6000 16.4000 113.8000 ;
	    RECT 15.4000 113.3000 16.4000 113.6000 ;
	    RECT 16.7000 113.4000 17.1000 113.5000 ;
	    RECT 15.4000 113.2000 16.2000 113.3000 ;
	    RECT 16.7000 113.1000 17.8000 113.4000 ;
	    RECT 14.8000 111.1000 15.6000 112.9000 ;
	    RECT 17.4000 111.1000 17.8000 113.1000 ;
	    RECT 18.2000 112.4000 18.6000 113.2000 ;
	    RECT 19.0000 111.1000 19.4000 119.9000 ;
	    RECT 19.8000 116.2000 20.2000 119.9000 ;
	    RECT 19.8000 115.9000 20.9000 116.2000 ;
	    RECT 20.6000 115.6000 20.9000 115.9000 ;
	    RECT 22.2000 115.6000 22.6000 119.9000 ;
	    RECT 24.3000 117.9000 24.9000 119.9000 ;
	    RECT 26.6000 117.9000 27.0000 119.9000 ;
	    RECT 28.8000 118.2000 29.2000 119.9000 ;
	    RECT 28.8000 117.9000 29.8000 118.2000 ;
	    RECT 24.6000 117.5000 25.0000 117.9000 ;
	    RECT 26.7000 117.6000 27.0000 117.9000 ;
	    RECT 26.3000 117.3000 28.1000 117.6000 ;
	    RECT 29.4000 117.5000 29.8000 117.9000 ;
	    RECT 26.3000 117.2000 26.7000 117.3000 ;
	    RECT 27.7000 117.2000 28.1000 117.3000 ;
	    RECT 24.2000 116.6000 24.9000 117.0000 ;
	    RECT 24.6000 116.1000 24.9000 116.6000 ;
	    RECT 25.7000 116.5000 26.8000 116.8000 ;
	    RECT 25.7000 116.4000 26.1000 116.5000 ;
	    RECT 24.6000 115.8000 25.8000 116.1000 ;
	    RECT 20.6000 115.2000 21.2000 115.6000 ;
	    RECT 22.2000 115.3000 24.3000 115.6000 ;
	    RECT 19.8000 114.4000 20.2000 115.2000 ;
	    RECT 20.6000 113.7000 20.9000 115.2000 ;
	    RECT 19.8000 113.4000 20.9000 113.7000 ;
	    RECT 22.2000 113.6000 22.6000 115.3000 ;
	    RECT 23.9000 115.2000 24.3000 115.3000 ;
	    RECT 25.5000 115.2000 25.8000 115.8000 ;
	    RECT 26.5000 115.9000 26.8000 116.5000 ;
	    RECT 27.1000 116.5000 27.5000 116.6000 ;
	    RECT 29.4000 116.5000 29.8000 116.6000 ;
	    RECT 27.1000 116.2000 29.8000 116.5000 ;
	    RECT 26.5000 115.7000 28.9000 115.9000 ;
	    RECT 31.0000 115.7000 31.4000 119.9000 ;
	    RECT 31.8000 116.2000 32.2000 119.9000 ;
	    RECT 32.6000 116.2000 33.0000 116.3000 ;
	    RECT 31.8000 115.9000 33.0000 116.2000 ;
	    RECT 34.0000 115.9000 34.8000 119.9000 ;
	    RECT 35.7000 116.2000 36.1000 116.3000 ;
	    RECT 36.6000 116.2000 37.0000 119.9000 ;
	    RECT 35.7000 115.9000 37.0000 116.2000 ;
	    RECT 38.7000 116.2000 39.1000 119.9000 ;
	    RECT 39.4000 116.8000 39.8000 117.2000 ;
	    RECT 39.5000 116.2000 39.8000 116.8000 ;
	    RECT 40.6000 116.2000 41.0000 119.9000 ;
	    RECT 42.2000 116.2000 42.6000 119.9000 ;
	    RECT 38.7000 115.9000 39.2000 116.2000 ;
	    RECT 39.5000 115.9000 40.2000 116.2000 ;
	    RECT 40.6000 115.9000 42.6000 116.2000 ;
	    RECT 43.0000 115.9000 43.4000 119.9000 ;
	    RECT 44.1000 116.3000 44.5000 119.9000 ;
	    RECT 44.1000 115.9000 45.0000 116.3000 ;
	    RECT 46.2000 116.2000 46.6000 119.9000 ;
	    RECT 50.3000 119.6000 52.1000 119.9000 ;
	    RECT 50.3000 119.5000 50.6000 119.6000 ;
	    RECT 50.2000 116.5000 50.6000 119.5000 ;
	    RECT 51.8000 119.5000 52.1000 119.6000 ;
	    RECT 52.6000 119.6000 54.6000 119.9000 ;
	    RECT 51.0000 116.5000 51.4000 119.3000 ;
	    RECT 51.8000 116.7000 52.2000 119.5000 ;
	    RECT 52.6000 117.0000 53.0000 119.6000 ;
	    RECT 53.4000 116.9000 53.8000 119.3000 ;
	    RECT 54.2000 116.9000 54.6000 119.6000 ;
	    RECT 53.4000 116.7000 53.7000 116.9000 ;
	    RECT 51.8000 116.5000 53.7000 116.7000 ;
	    RECT 51.1000 116.2000 51.4000 116.5000 ;
	    RECT 51.9000 116.4000 53.7000 116.5000 ;
	    RECT 54.3000 116.6000 54.6000 116.9000 ;
	    RECT 55.8000 116.9000 56.2000 119.9000 ;
	    RECT 55.8000 116.6000 56.1000 116.9000 ;
	    RECT 54.3000 116.3000 56.1000 116.6000 ;
	    RECT 56.9000 116.3000 57.3000 119.9000 ;
	    RECT 46.2000 115.9000 47.3000 116.2000 ;
	    RECT 26.5000 115.6000 31.4000 115.7000 ;
	    RECT 28.5000 115.5000 31.4000 115.6000 ;
	    RECT 28.6000 115.4000 31.4000 115.5000 ;
	    RECT 34.2000 115.2000 34.5000 115.9000 ;
	    RECT 35.1000 115.2000 35.5000 115.3000 ;
	    RECT 23.1000 114.9000 23.5000 115.0000 ;
	    RECT 23.1000 114.6000 25.0000 114.9000 ;
	    RECT 25.4000 114.8000 25.8000 115.2000 ;
	    RECT 27.8000 115.1000 28.2000 115.2000 ;
	    RECT 27.8000 114.8000 30.3000 115.1000 ;
	    RECT 24.6000 114.5000 25.0000 114.6000 ;
	    RECT 25.5000 114.2000 25.8000 114.8000 ;
	    RECT 28.6000 114.7000 29.0000 114.8000 ;
	    RECT 29.9000 114.7000 30.3000 114.8000 ;
	    RECT 34.2000 114.8000 34.6000 115.2000 ;
	    RECT 35.1000 114.9000 35.9000 115.2000 ;
	    RECT 35.5000 114.8000 35.9000 114.9000 ;
	    RECT 29.1000 114.2000 29.5000 114.3000 ;
	    RECT 34.2000 114.2000 34.5000 114.8000 ;
	    RECT 38.2000 114.4000 38.6000 115.2000 ;
	    RECT 38.9000 115.1000 39.2000 115.9000 ;
	    RECT 39.8000 115.8000 40.2000 115.9000 ;
	    RECT 41.0000 115.2000 41.4000 115.4000 ;
	    RECT 43.0000 115.2000 43.3000 115.9000 ;
	    RECT 39.8000 115.1000 40.2000 115.2000 ;
	    RECT 38.9000 114.8000 40.2000 115.1000 ;
	    RECT 40.6000 114.9000 41.4000 115.2000 ;
	    RECT 42.2000 115.1000 43.4000 115.2000 ;
	    RECT 43.8000 115.1000 44.2000 115.6000 ;
	    RECT 42.2000 114.9000 44.2000 115.1000 ;
	    RECT 40.6000 114.8000 41.0000 114.9000 ;
	    RECT 25.5000 113.9000 31.0000 114.2000 ;
	    RECT 25.7000 113.8000 26.1000 113.9000 ;
	    RECT 19.8000 111.1000 20.2000 113.4000 ;
	    RECT 22.2000 113.3000 24.1000 113.6000 ;
	    RECT 22.2000 111.1000 22.6000 113.3000 ;
	    RECT 23.7000 113.2000 24.1000 113.3000 ;
	    RECT 28.6000 112.8000 28.9000 113.9000 ;
	    RECT 30.2000 113.8000 31.0000 113.9000 ;
	    RECT 31.8000 113.8000 32.6000 114.2000 ;
	    RECT 33.2000 113.8000 33.6000 114.2000 ;
	    RECT 33.3000 113.6000 33.6000 113.8000 ;
	    RECT 34.0000 113.9000 34.5000 114.2000 ;
	    RECT 34.8000 114.3000 35.2000 114.4000 ;
	    RECT 34.8000 114.2000 36.2000 114.3000 ;
	    RECT 38.9000 114.2000 39.2000 114.8000 ;
	    RECT 34.8000 114.0000 37.0000 114.2000 ;
	    RECT 35.9000 113.9000 37.0000 114.0000 ;
	    RECT 27.7000 112.7000 28.1000 112.8000 ;
	    RECT 24.6000 112.1000 25.0000 112.5000 ;
	    RECT 26.7000 112.4000 28.1000 112.7000 ;
	    RECT 28.6000 112.4000 29.0000 112.8000 ;
	    RECT 26.7000 112.1000 27.0000 112.4000 ;
	    RECT 29.4000 112.1000 29.8000 112.5000 ;
	    RECT 24.3000 111.8000 25.0000 112.1000 ;
	    RECT 24.3000 111.1000 24.9000 111.8000 ;
	    RECT 26.6000 111.1000 27.0000 112.1000 ;
	    RECT 28.8000 111.8000 29.8000 112.1000 ;
	    RECT 28.8000 111.1000 29.2000 111.8000 ;
	    RECT 31.0000 111.1000 31.4000 113.5000 ;
	    RECT 32.6000 113.4000 33.0000 113.5000 ;
	    RECT 31.8000 113.1000 33.0000 113.4000 ;
	    RECT 33.3000 113.2000 33.7000 113.6000 ;
	    RECT 31.8000 111.1000 32.2000 113.1000 ;
	    RECT 34.0000 112.9000 34.3000 113.9000 ;
	    RECT 36.2000 113.8000 37.0000 113.9000 ;
	    RECT 37.4000 114.1000 37.8000 114.2000 ;
	    RECT 37.4000 113.8000 38.2000 114.1000 ;
	    RECT 38.9000 113.8000 40.2000 114.2000 ;
	    RECT 41.4000 113.8000 41.8000 114.6000 ;
	    RECT 37.8000 113.6000 38.2000 113.8000 ;
	    RECT 34.6000 113.2000 35.4000 113.6000 ;
	    RECT 35.7000 113.4000 36.1000 113.5000 ;
	    RECT 35.7000 113.1000 37.0000 113.4000 ;
	    RECT 37.5000 113.1000 39.3000 113.3000 ;
	    RECT 39.8000 113.1000 40.1000 113.8000 ;
	    RECT 42.2000 113.1000 42.5000 114.9000 ;
	    RECT 43.0000 114.8000 44.2000 114.9000 ;
	    RECT 43.8000 114.2000 44.1000 114.8000 ;
	    RECT 44.6000 114.2000 44.9000 115.9000 ;
	    RECT 47.0000 115.6000 47.3000 115.9000 ;
	    RECT 51.0000 116.1000 51.4000 116.2000 ;
	    RECT 51.0000 115.8000 52.7000 116.1000 ;
	    RECT 56.9000 115.9000 57.8000 116.3000 ;
	    RECT 59.0000 116.2000 59.4000 119.9000 ;
	    RECT 59.7000 116.2000 60.1000 116.3000 ;
	    RECT 59.0000 115.9000 60.1000 116.2000 ;
	    RECT 61.2000 116.2000 62.0000 119.9000 ;
	    RECT 63.0000 116.2000 63.4000 116.3000 ;
	    RECT 63.8000 116.2000 64.2000 119.9000 ;
	    RECT 61.2000 115.9000 62.2000 116.2000 ;
	    RECT 63.0000 115.9000 64.2000 116.2000 ;
	    RECT 47.0000 115.2000 47.6000 115.6000 ;
	    RECT 46.2000 114.4000 46.6000 115.2000 ;
	    RECT 43.8000 113.8000 44.2000 114.2000 ;
	    RECT 44.6000 113.8000 45.0000 114.2000 ;
	    RECT 34.0000 112.2000 34.8000 112.9000 ;
	    RECT 33.4000 111.8000 34.8000 112.2000 ;
	    RECT 34.0000 111.1000 34.8000 111.8000 ;
	    RECT 36.6000 111.1000 37.0000 113.1000 ;
	    RECT 37.4000 113.0000 39.4000 113.1000 ;
	    RECT 37.4000 111.1000 37.8000 113.0000 ;
	    RECT 39.0000 111.1000 39.4000 113.0000 ;
	    RECT 39.8000 111.1000 40.2000 113.1000 ;
	    RECT 42.2000 111.1000 42.6000 113.1000 ;
	    RECT 43.0000 112.8000 43.4000 113.2000 ;
	    RECT 43.8000 113.1000 44.2000 113.2000 ;
	    RECT 44.6000 113.1000 44.9000 113.8000 ;
	    RECT 47.0000 113.7000 47.3000 115.2000 ;
	    RECT 46.2000 113.4000 47.3000 113.7000 ;
	    RECT 43.8000 112.8000 44.9000 113.1000 ;
	    RECT 42.9000 112.4000 43.3000 112.8000 ;
	    RECT 44.6000 112.1000 44.9000 112.8000 ;
	    RECT 45.4000 112.4000 45.8000 113.2000 ;
	    RECT 44.6000 111.1000 45.0000 112.1000 ;
	    RECT 46.2000 111.1000 46.6000 113.4000 ;
	    RECT 52.4000 112.5000 52.7000 115.8000 ;
	    RECT 53.0000 115.1000 53.8000 115.2000 ;
	    RECT 56.6000 115.1000 57.0000 115.6000 ;
	    RECT 53.0000 114.8000 57.0000 115.1000 ;
	    RECT 57.4000 114.2000 57.7000 115.9000 ;
	    RECT 59.8000 115.6000 60.1000 115.9000 ;
	    RECT 59.8000 115.3000 61.5000 115.6000 ;
	    RECT 61.1000 115.2000 61.5000 115.3000 ;
	    RECT 61.9000 115.2000 62.2000 115.9000 ;
	    RECT 64.6000 115.8000 65.0000 116.6000 ;
	    RECT 61.9000 115.1000 62.6000 115.2000 ;
	    RECT 63.8000 115.1000 64.2000 115.2000 ;
	    RECT 60.0000 114.9000 60.4000 115.0000 ;
	    RECT 61.9000 114.9000 64.2000 115.1000 ;
	    RECT 60.0000 114.6000 61.3000 114.9000 ;
	    RECT 61.0000 114.3000 61.3000 114.6000 ;
	    RECT 61.7000 114.8000 64.2000 114.9000 ;
	    RECT 61.7000 114.6000 62.2000 114.8000 ;
	    RECT 53.8000 113.8000 54.6000 114.2000 ;
	    RECT 57.4000 114.1000 57.8000 114.2000 ;
	    RECT 59.0000 114.1000 59.8000 114.2000 ;
	    RECT 57.4000 113.8000 60.7000 114.1000 ;
	    RECT 61.0000 113.9000 61.4000 114.3000 ;
	    RECT 54.5000 112.8000 55.4000 113.2000 ;
	    RECT 52.4000 112.2000 54.4000 112.5000 ;
	    RECT 52.4000 112.1000 53.0000 112.2000 ;
	    RECT 52.6000 111.1000 53.0000 112.1000 ;
	    RECT 54.1000 112.1000 54.4000 112.2000 ;
	    RECT 57.4000 112.1000 57.7000 113.8000 ;
	    RECT 60.4000 113.6000 60.7000 113.8000 ;
	    RECT 59.7000 113.4000 60.1000 113.5000 ;
	    RECT 58.2000 112.4000 58.6000 113.2000 ;
	    RECT 59.0000 113.1000 60.1000 113.4000 ;
	    RECT 60.4000 113.3000 61.4000 113.6000 ;
	    RECT 60.6000 113.2000 61.4000 113.3000 ;
	    RECT 54.1000 111.8000 54.6000 112.1000 ;
	    RECT 54.2000 111.1000 54.6000 111.8000 ;
	    RECT 57.4000 111.1000 57.8000 112.1000 ;
	    RECT 59.0000 111.1000 59.4000 113.1000 ;
	    RECT 61.7000 112.9000 62.0000 114.6000 ;
	    RECT 62.4000 113.8000 62.8000 114.2000 ;
	    RECT 63.4000 114.1000 64.2000 114.2000 ;
	    RECT 64.6000 114.1000 65.0000 114.2000 ;
	    RECT 63.4000 113.8000 65.0000 114.1000 ;
	    RECT 62.4000 113.6000 62.7000 113.8000 ;
	    RECT 62.3000 113.2000 62.7000 113.6000 ;
	    RECT 63.0000 113.4000 63.4000 113.5000 ;
	    RECT 63.0000 113.1000 64.2000 113.4000 ;
	    RECT 65.4000 113.1000 65.8000 119.9000 ;
	    RECT 66.2000 116.8000 66.6000 117.2000 ;
	    RECT 66.2000 116.1000 66.5000 116.8000 ;
	    RECT 67.0000 116.1000 67.4000 119.9000 ;
	    RECT 66.2000 115.8000 67.4000 116.1000 ;
	    RECT 68.6000 116.2000 69.0000 119.9000 ;
	    RECT 68.6000 115.9000 69.7000 116.2000 ;
	    RECT 66.2000 113.4000 66.6000 114.2000 ;
	    RECT 61.2000 111.1000 62.0000 112.9000 ;
	    RECT 63.8000 111.1000 64.2000 113.1000 ;
	    RECT 64.9000 112.8000 65.8000 113.1000 ;
	    RECT 64.9000 112.2000 65.3000 112.8000 ;
	    RECT 64.6000 111.8000 65.3000 112.2000 ;
	    RECT 64.9000 111.1000 65.3000 111.8000 ;
	    RECT 67.0000 111.1000 67.4000 115.8000 ;
	    RECT 69.4000 115.6000 69.7000 115.9000 ;
	    RECT 71.0000 115.7000 71.4000 119.9000 ;
	    RECT 73.2000 118.2000 73.6000 119.9000 ;
	    RECT 72.6000 117.9000 73.6000 118.2000 ;
	    RECT 75.4000 117.9000 75.8000 119.9000 ;
	    RECT 77.5000 117.9000 78.1000 119.9000 ;
	    RECT 72.6000 117.5000 73.0000 117.9000 ;
	    RECT 75.4000 117.6000 75.7000 117.9000 ;
	    RECT 74.3000 117.3000 76.1000 117.6000 ;
	    RECT 77.4000 117.5000 77.8000 117.9000 ;
	    RECT 74.3000 117.2000 74.7000 117.3000 ;
	    RECT 75.7000 117.2000 76.1000 117.3000 ;
	    RECT 72.6000 116.5000 73.0000 116.6000 ;
	    RECT 74.9000 116.5000 75.3000 116.6000 ;
	    RECT 72.6000 116.2000 75.3000 116.5000 ;
	    RECT 75.6000 116.5000 76.7000 116.8000 ;
	    RECT 75.6000 115.9000 75.9000 116.5000 ;
	    RECT 76.3000 116.4000 76.7000 116.5000 ;
	    RECT 77.5000 116.6000 78.2000 117.0000 ;
	    RECT 77.5000 116.1000 77.8000 116.6000 ;
	    RECT 73.5000 115.7000 75.9000 115.9000 ;
	    RECT 71.0000 115.6000 75.9000 115.7000 ;
	    RECT 76.6000 115.8000 77.8000 116.1000 ;
	    RECT 69.4000 115.2000 70.0000 115.6000 ;
	    RECT 71.0000 115.5000 73.9000 115.6000 ;
	    RECT 71.0000 115.4000 73.8000 115.5000 ;
	    RECT 68.6000 114.4000 69.0000 115.2000 ;
	    RECT 67.8000 113.4000 68.2000 114.2000 ;
	    RECT 69.4000 113.7000 69.7000 115.2000 ;
	    RECT 74.2000 115.1000 74.6000 115.2000 ;
	    RECT 72.1000 114.8000 74.6000 115.1000 ;
	    RECT 72.1000 114.7000 72.5000 114.8000 ;
	    RECT 73.4000 114.7000 73.8000 114.8000 ;
	    RECT 72.9000 114.2000 73.3000 114.3000 ;
	    RECT 76.6000 114.2000 76.9000 115.8000 ;
	    RECT 79.8000 115.6000 80.2000 119.9000 ;
	    RECT 80.6000 116.2000 81.0000 119.9000 ;
	    RECT 83.0000 116.2000 83.4000 119.9000 ;
	    RECT 85.4000 116.2000 85.8000 119.9000 ;
	    RECT 87.8000 116.2000 88.2000 119.9000 ;
	    RECT 90.2000 116.2000 90.6000 119.9000 ;
	    RECT 92.6000 116.2000 93.0000 119.9000 ;
	    RECT 95.0000 116.2000 95.4000 119.9000 ;
	    RECT 95.9000 116.2000 96.3000 116.3000 ;
	    RECT 80.6000 115.9000 81.7000 116.2000 ;
	    RECT 83.0000 115.9000 84.1000 116.2000 ;
	    RECT 85.4000 115.9000 86.5000 116.2000 ;
	    RECT 87.8000 115.9000 88.9000 116.2000 ;
	    RECT 90.2000 115.9000 91.3000 116.2000 ;
	    RECT 92.6000 115.9000 93.7000 116.2000 ;
	    RECT 95.0000 115.9000 96.3000 116.2000 ;
	    RECT 97.2000 115.9000 98.0000 119.9000 ;
	    RECT 99.0000 116.2000 99.4000 116.3000 ;
	    RECT 99.8000 116.2000 100.2000 119.9000 ;
	    RECT 99.0000 115.9000 100.2000 116.2000 ;
	    RECT 102.2000 116.2000 102.6000 119.9000 ;
	    RECT 104.6000 116.2000 105.0000 119.9000 ;
	    RECT 102.2000 115.9000 103.3000 116.2000 ;
	    RECT 104.6000 115.9000 105.7000 116.2000 ;
	    RECT 78.1000 115.3000 80.2000 115.6000 ;
	    RECT 78.1000 115.2000 78.5000 115.3000 ;
	    RECT 79.8000 115.1000 80.2000 115.3000 ;
	    RECT 81.4000 115.6000 81.7000 115.9000 ;
	    RECT 83.8000 115.6000 84.1000 115.9000 ;
	    RECT 86.2000 115.6000 86.5000 115.9000 ;
	    RECT 88.6000 115.6000 88.9000 115.9000 ;
	    RECT 91.0000 115.6000 91.3000 115.9000 ;
	    RECT 93.4000 115.6000 93.7000 115.9000 ;
	    RECT 81.4000 115.2000 82.0000 115.6000 ;
	    RECT 83.8000 115.2000 84.4000 115.6000 ;
	    RECT 86.2000 115.2000 86.8000 115.6000 ;
	    RECT 88.6000 115.2000 89.2000 115.6000 ;
	    RECT 91.0000 115.2000 91.6000 115.6000 ;
	    RECT 93.4000 115.2000 94.0000 115.6000 ;
	    RECT 96.5000 115.2000 96.9000 115.3000 ;
	    RECT 97.5000 115.2000 97.8000 115.9000 ;
	    RECT 103.0000 115.6000 103.3000 115.9000 ;
	    RECT 105.4000 115.6000 105.7000 115.9000 ;
	    RECT 103.0000 115.2000 103.6000 115.6000 ;
	    RECT 105.4000 115.2000 106.0000 115.6000 ;
	    RECT 80.6000 115.1000 81.0000 115.2000 ;
	    RECT 78.9000 114.9000 79.3000 115.0000 ;
	    RECT 77.4000 114.6000 79.3000 114.9000 ;
	    RECT 79.8000 114.8000 81.0000 115.1000 ;
	    RECT 77.4000 114.5000 77.8000 114.6000 ;
	    RECT 71.4000 113.9000 76.9000 114.2000 ;
	    RECT 71.4000 113.8000 72.2000 113.9000 ;
	    RECT 68.6000 113.4000 69.7000 113.7000 ;
	    RECT 68.6000 111.1000 69.0000 113.4000 ;
	    RECT 71.0000 111.1000 71.4000 113.5000 ;
	    RECT 73.5000 112.8000 73.8000 113.9000 ;
	    RECT 75.0000 113.8000 75.4000 113.9000 ;
	    RECT 76.3000 113.8000 76.7000 113.9000 ;
	    RECT 78.2000 113.6000 78.6000 114.2000 ;
	    RECT 79.8000 113.6000 80.2000 114.8000 ;
	    RECT 80.6000 114.4000 81.0000 114.8000 ;
	    RECT 81.4000 113.7000 81.7000 115.2000 ;
	    RECT 83.0000 114.4000 83.4000 115.2000 ;
	    RECT 83.8000 113.7000 84.1000 115.2000 ;
	    RECT 85.4000 114.4000 85.8000 115.2000 ;
	    RECT 86.2000 113.7000 86.5000 115.2000 ;
	    RECT 87.8000 114.4000 88.2000 115.2000 ;
	    RECT 88.6000 113.7000 88.9000 115.2000 ;
	    RECT 90.2000 114.4000 90.6000 115.2000 ;
	    RECT 91.0000 113.7000 91.3000 115.2000 ;
	    RECT 92.6000 114.4000 93.0000 115.2000 ;
	    RECT 93.4000 113.7000 93.7000 115.2000 ;
	    RECT 96.1000 114.9000 96.9000 115.2000 ;
	    RECT 96.1000 114.8000 96.5000 114.9000 ;
	    RECT 97.4000 114.8000 97.8000 115.2000 ;
	    RECT 102.2000 115.1000 102.6000 115.2000 ;
	    RECT 96.8000 114.3000 97.2000 114.4000 ;
	    RECT 95.8000 114.2000 97.2000 114.3000 ;
	    RECT 95.0000 114.0000 97.2000 114.2000 ;
	    RECT 97.5000 114.2000 97.8000 114.8000 ;
	    RECT 99.8000 114.8000 102.6000 115.1000 ;
	    RECT 99.8000 114.2000 100.1000 114.8000 ;
	    RECT 102.2000 114.4000 102.6000 114.8000 ;
	    RECT 95.0000 113.9000 96.1000 114.0000 ;
	    RECT 97.5000 113.9000 98.0000 114.2000 ;
	    RECT 95.0000 113.8000 95.8000 113.9000 ;
	    RECT 78.2000 113.3000 80.2000 113.6000 ;
	    RECT 78.3000 113.2000 78.7000 113.3000 ;
	    RECT 72.6000 112.1000 73.0000 112.5000 ;
	    RECT 73.4000 112.4000 73.8000 112.8000 ;
	    RECT 74.3000 112.7000 74.7000 112.8000 ;
	    RECT 74.3000 112.4000 75.7000 112.7000 ;
	    RECT 75.4000 112.1000 75.7000 112.4000 ;
	    RECT 77.4000 112.1000 77.8000 112.5000 ;
	    RECT 72.6000 111.8000 73.6000 112.1000 ;
	    RECT 73.2000 111.1000 73.6000 111.8000 ;
	    RECT 75.4000 111.1000 75.8000 112.1000 ;
	    RECT 77.4000 111.8000 78.1000 112.1000 ;
	    RECT 77.5000 111.1000 78.1000 111.8000 ;
	    RECT 79.8000 111.1000 80.2000 113.3000 ;
	    RECT 80.6000 113.4000 81.7000 113.7000 ;
	    RECT 83.0000 113.4000 84.1000 113.7000 ;
	    RECT 85.4000 113.4000 86.5000 113.7000 ;
	    RECT 87.8000 113.4000 88.9000 113.7000 ;
	    RECT 90.2000 113.4000 91.3000 113.7000 ;
	    RECT 92.6000 113.4000 93.7000 113.7000 ;
	    RECT 95.9000 113.4000 96.3000 113.5000 ;
	    RECT 80.6000 111.1000 81.0000 113.4000 ;
	    RECT 83.0000 111.1000 83.4000 113.4000 ;
	    RECT 85.4000 111.1000 85.8000 113.4000 ;
	    RECT 87.8000 111.1000 88.2000 113.4000 ;
	    RECT 90.2000 111.1000 90.6000 113.4000 ;
	    RECT 92.6000 111.1000 93.0000 113.4000 ;
	    RECT 95.0000 113.1000 96.3000 113.4000 ;
	    RECT 96.6000 113.2000 97.4000 113.6000 ;
	    RECT 95.0000 111.1000 95.4000 113.1000 ;
	    RECT 97.7000 112.9000 98.0000 113.9000 ;
	    RECT 98.4000 113.8000 98.8000 114.2000 ;
	    RECT 99.4000 113.8000 100.2000 114.2000 ;
	    RECT 98.4000 113.6000 98.7000 113.8000 ;
	    RECT 103.0000 113.7000 103.3000 115.2000 ;
	    RECT 104.6000 114.4000 105.0000 115.2000 ;
	    RECT 105.4000 113.7000 105.7000 115.2000 ;
	    RECT 98.3000 113.2000 98.7000 113.6000 ;
	    RECT 99.0000 113.4000 99.4000 113.5000 ;
	    RECT 102.2000 113.4000 103.3000 113.7000 ;
	    RECT 104.6000 113.4000 105.7000 113.7000 ;
	    RECT 107.0000 113.4000 107.4000 114.2000 ;
	    RECT 99.0000 113.1000 100.2000 113.4000 ;
	    RECT 97.2000 112.2000 98.0000 112.9000 ;
	    RECT 97.2000 111.8000 98.6000 112.2000 ;
	    RECT 97.2000 111.1000 98.0000 111.8000 ;
	    RECT 99.8000 111.1000 100.2000 113.1000 ;
	    RECT 102.2000 111.1000 102.6000 113.4000 ;
	    RECT 104.6000 111.1000 105.0000 113.4000 ;
	    RECT 107.8000 113.1000 108.2000 119.9000 ;
	    RECT 109.4000 113.4000 109.8000 114.2000 ;
	    RECT 110.2000 113.1000 110.6000 119.9000 ;
	    RECT 111.8000 115.7000 112.2000 119.9000 ;
	    RECT 114.0000 118.2000 114.4000 119.9000 ;
	    RECT 113.4000 117.9000 114.4000 118.2000 ;
	    RECT 116.2000 117.9000 116.6000 119.9000 ;
	    RECT 118.3000 117.9000 118.9000 119.9000 ;
	    RECT 113.4000 117.5000 113.8000 117.9000 ;
	    RECT 116.2000 117.6000 116.5000 117.9000 ;
	    RECT 115.1000 117.3000 116.9000 117.6000 ;
	    RECT 118.2000 117.5000 118.6000 117.9000 ;
	    RECT 115.1000 117.2000 115.5000 117.3000 ;
	    RECT 116.5000 117.2000 116.9000 117.3000 ;
	    RECT 113.4000 116.5000 113.8000 116.6000 ;
	    RECT 115.7000 116.5000 116.1000 116.6000 ;
	    RECT 113.4000 116.2000 116.1000 116.5000 ;
	    RECT 116.4000 116.5000 117.5000 116.8000 ;
	    RECT 116.4000 115.9000 116.7000 116.5000 ;
	    RECT 117.1000 116.4000 117.5000 116.5000 ;
	    RECT 118.3000 116.6000 119.0000 117.0000 ;
	    RECT 118.3000 116.1000 118.6000 116.6000 ;
	    RECT 114.3000 115.7000 116.7000 115.9000 ;
	    RECT 111.8000 115.6000 116.7000 115.7000 ;
	    RECT 117.4000 115.8000 118.6000 116.1000 ;
	    RECT 111.8000 115.5000 114.7000 115.6000 ;
	    RECT 111.8000 115.4000 114.6000 115.5000 ;
	    RECT 115.0000 115.1000 115.4000 115.2000 ;
	    RECT 112.9000 114.8000 115.4000 115.1000 ;
	    RECT 116.6000 115.1000 117.0000 115.2000 ;
	    RECT 117.4000 115.1000 117.7000 115.8000 ;
	    RECT 120.6000 115.6000 121.0000 119.9000 ;
	    RECT 121.4000 116.2000 121.8000 119.9000 ;
	    RECT 125.4000 116.2000 125.8000 119.9000 ;
	    RECT 121.4000 115.9000 122.5000 116.2000 ;
	    RECT 118.9000 115.3000 121.0000 115.6000 ;
	    RECT 118.9000 115.2000 119.3000 115.3000 ;
	    RECT 116.6000 114.8000 117.7000 115.1000 ;
	    RECT 120.6000 115.1000 121.0000 115.3000 ;
	    RECT 122.2000 115.6000 122.5000 115.9000 ;
	    RECT 124.7000 115.9000 125.8000 116.2000 ;
	    RECT 124.7000 115.6000 125.0000 115.9000 ;
	    RECT 122.2000 115.2000 122.8000 115.6000 ;
	    RECT 124.4000 115.2000 125.0000 115.6000 ;
	    RECT 126.2000 115.6000 126.6000 119.9000 ;
	    RECT 128.3000 117.9000 128.9000 119.9000 ;
	    RECT 130.6000 117.9000 131.0000 119.9000 ;
	    RECT 132.8000 118.2000 133.2000 119.9000 ;
	    RECT 132.8000 117.9000 133.8000 118.2000 ;
	    RECT 128.6000 117.5000 129.0000 117.9000 ;
	    RECT 130.7000 117.6000 131.0000 117.9000 ;
	    RECT 130.3000 117.3000 132.1000 117.6000 ;
	    RECT 133.4000 117.5000 133.8000 117.9000 ;
	    RECT 130.3000 117.2000 130.7000 117.3000 ;
	    RECT 131.7000 117.2000 132.1000 117.3000 ;
	    RECT 128.2000 116.6000 128.9000 117.0000 ;
	    RECT 128.6000 116.1000 128.9000 116.6000 ;
	    RECT 129.7000 116.5000 130.8000 116.8000 ;
	    RECT 129.7000 116.4000 130.1000 116.5000 ;
	    RECT 128.6000 115.8000 129.8000 116.1000 ;
	    RECT 126.2000 115.3000 128.3000 115.6000 ;
	    RECT 121.4000 115.1000 121.8000 115.2000 ;
	    RECT 119.7000 114.9000 120.1000 115.0000 ;
	    RECT 112.9000 114.7000 113.3000 114.8000 ;
	    RECT 113.7000 114.2000 114.1000 114.3000 ;
	    RECT 117.4000 114.2000 117.7000 114.8000 ;
	    RECT 118.2000 114.6000 120.1000 114.9000 ;
	    RECT 120.6000 114.8000 121.8000 115.1000 ;
	    RECT 118.2000 114.5000 118.6000 114.6000 ;
	    RECT 112.2000 113.9000 117.7000 114.2000 ;
	    RECT 112.2000 113.8000 113.0000 113.9000 ;
	    RECT 107.8000 112.8000 108.7000 113.1000 ;
	    RECT 110.2000 112.8000 111.1000 113.1000 ;
	    RECT 108.3000 112.2000 108.7000 112.8000 ;
	    RECT 110.7000 112.2000 111.1000 112.8000 ;
	    RECT 108.3000 111.8000 109.0000 112.2000 ;
	    RECT 110.7000 111.8000 111.4000 112.2000 ;
	    RECT 108.3000 111.1000 108.7000 111.8000 ;
	    RECT 110.7000 111.1000 111.1000 111.8000 ;
	    RECT 111.8000 111.1000 112.2000 113.5000 ;
	    RECT 114.3000 112.8000 114.6000 113.9000 ;
	    RECT 117.1000 113.8000 117.5000 113.9000 ;
	    RECT 120.6000 113.6000 121.0000 114.8000 ;
	    RECT 121.4000 114.4000 121.8000 114.8000 ;
	    RECT 122.2000 113.7000 122.5000 115.2000 ;
	    RECT 119.1000 113.3000 121.0000 113.6000 ;
	    RECT 119.1000 113.2000 119.5000 113.3000 ;
	    RECT 113.4000 112.1000 113.8000 112.5000 ;
	    RECT 114.2000 112.4000 114.6000 112.8000 ;
	    RECT 115.1000 112.7000 115.5000 112.8000 ;
	    RECT 115.1000 112.4000 116.5000 112.7000 ;
	    RECT 116.2000 112.1000 116.5000 112.4000 ;
	    RECT 118.2000 112.1000 118.6000 112.5000 ;
	    RECT 113.4000 111.8000 114.4000 112.1000 ;
	    RECT 114.0000 111.1000 114.4000 111.8000 ;
	    RECT 116.2000 111.1000 116.6000 112.1000 ;
	    RECT 118.2000 111.8000 118.9000 112.1000 ;
	    RECT 118.3000 111.1000 118.9000 111.8000 ;
	    RECT 120.6000 111.1000 121.0000 113.3000 ;
	    RECT 121.4000 113.4000 122.5000 113.7000 ;
	    RECT 124.7000 113.7000 125.0000 115.2000 ;
	    RECT 125.4000 115.1000 125.8000 115.2000 ;
	    RECT 126.2000 115.1000 126.6000 115.3000 ;
	    RECT 127.9000 115.2000 128.3000 115.3000 ;
	    RECT 129.5000 115.2000 129.8000 115.8000 ;
	    RECT 130.5000 115.9000 130.8000 116.5000 ;
	    RECT 131.1000 116.5000 131.5000 116.6000 ;
	    RECT 133.4000 116.5000 133.8000 116.6000 ;
	    RECT 131.1000 116.2000 133.8000 116.5000 ;
	    RECT 130.5000 115.7000 132.9000 115.9000 ;
	    RECT 135.0000 115.7000 135.4000 119.9000 ;
	    RECT 135.8000 116.2000 136.2000 119.9000 ;
	    RECT 135.8000 115.9000 136.9000 116.2000 ;
	    RECT 130.5000 115.6000 135.4000 115.7000 ;
	    RECT 132.5000 115.5000 135.4000 115.6000 ;
	    RECT 132.6000 115.4000 135.4000 115.5000 ;
	    RECT 136.6000 115.6000 136.9000 115.9000 ;
	    RECT 138.2000 115.9000 138.6000 119.9000 ;
	    RECT 139.8000 116.2000 140.2000 119.9000 ;
	    RECT 139.1000 115.9000 140.2000 116.2000 ;
	    RECT 140.6000 116.2000 141.0000 119.9000 ;
	    RECT 143.0000 116.2000 143.4000 119.9000 ;
	    RECT 145.4000 116.2000 145.8000 119.9000 ;
	    RECT 140.6000 115.9000 141.7000 116.2000 ;
	    RECT 143.0000 115.9000 144.1000 116.2000 ;
	    RECT 145.4000 115.9000 146.5000 116.2000 ;
	    RECT 136.6000 115.2000 137.2000 115.6000 ;
	    RECT 125.4000 114.8000 126.6000 115.1000 ;
	    RECT 125.4000 114.4000 125.8000 114.8000 ;
	    RECT 124.7000 113.4000 125.8000 113.7000 ;
	    RECT 121.4000 111.1000 121.8000 113.4000 ;
	    RECT 125.4000 111.1000 125.8000 113.4000 ;
	    RECT 126.2000 113.6000 126.6000 114.8000 ;
	    RECT 127.1000 114.9000 127.5000 115.0000 ;
	    RECT 127.1000 114.6000 129.0000 114.9000 ;
	    RECT 129.4000 114.8000 129.8000 115.2000 ;
	    RECT 131.8000 115.1000 132.2000 115.2000 ;
	    RECT 131.8000 114.8000 134.3000 115.1000 ;
	    RECT 128.6000 114.5000 129.0000 114.6000 ;
	    RECT 129.5000 114.2000 129.8000 114.8000 ;
	    RECT 132.6000 114.7000 133.0000 114.8000 ;
	    RECT 133.9000 114.7000 134.3000 114.8000 ;
	    RECT 135.8000 114.4000 136.2000 115.2000 ;
	    RECT 133.1000 114.2000 133.5000 114.3000 ;
	    RECT 129.5000 113.9000 135.0000 114.2000 ;
	    RECT 129.7000 113.8000 130.1000 113.9000 ;
	    RECT 126.2000 113.3000 128.2000 113.6000 ;
	    RECT 126.2000 111.1000 126.6000 113.3000 ;
	    RECT 127.7000 113.2000 128.2000 113.3000 ;
	    RECT 127.8000 113.1000 128.2000 113.2000 ;
	    RECT 129.4000 113.1000 129.8000 113.2000 ;
	    RECT 127.8000 112.8000 129.8000 113.1000 ;
	    RECT 132.6000 112.8000 132.9000 113.9000 ;
	    RECT 134.2000 113.8000 135.0000 113.9000 ;
	    RECT 136.6000 113.7000 136.9000 115.2000 ;
	    RECT 131.7000 112.7000 132.1000 112.8000 ;
	    RECT 128.6000 112.1000 129.0000 112.5000 ;
	    RECT 130.7000 112.4000 132.1000 112.7000 ;
	    RECT 132.6000 112.4000 133.0000 112.8000 ;
	    RECT 130.7000 112.1000 131.0000 112.4000 ;
	    RECT 133.4000 112.1000 133.8000 112.5000 ;
	    RECT 128.3000 111.8000 129.0000 112.1000 ;
	    RECT 128.3000 111.1000 128.9000 111.8000 ;
	    RECT 130.6000 111.1000 131.0000 112.1000 ;
	    RECT 132.8000 111.8000 133.8000 112.1000 ;
	    RECT 132.8000 111.1000 133.2000 111.8000 ;
	    RECT 135.0000 111.1000 135.4000 113.5000 ;
	    RECT 135.8000 113.4000 136.9000 113.7000 ;
	    RECT 138.2000 114.8000 138.5000 115.9000 ;
	    RECT 139.1000 115.6000 139.4000 115.9000 ;
	    RECT 138.8000 115.2000 139.4000 115.6000 ;
	    RECT 141.4000 115.6000 141.7000 115.9000 ;
	    RECT 143.8000 115.6000 144.1000 115.9000 ;
	    RECT 146.2000 115.6000 146.5000 115.9000 ;
	    RECT 141.4000 115.2000 142.0000 115.6000 ;
	    RECT 143.8000 115.2000 144.4000 115.6000 ;
	    RECT 146.2000 115.2000 146.8000 115.6000 ;
	    RECT 135.8000 111.1000 136.2000 113.4000 ;
	    RECT 138.2000 111.1000 138.6000 114.8000 ;
	    RECT 139.1000 113.7000 139.4000 115.2000 ;
	    RECT 139.8000 115.1000 140.2000 115.2000 ;
	    RECT 140.6000 115.1000 141.0000 115.2000 ;
	    RECT 139.8000 114.8000 141.0000 115.1000 ;
	    RECT 139.8000 114.4000 140.2000 114.8000 ;
	    RECT 140.6000 114.4000 141.0000 114.8000 ;
	    RECT 141.4000 113.7000 141.7000 115.2000 ;
	    RECT 143.0000 114.4000 143.4000 115.2000 ;
	    RECT 143.8000 113.7000 144.1000 115.2000 ;
	    RECT 145.4000 114.4000 145.8000 115.2000 ;
	    RECT 146.2000 113.7000 146.5000 115.2000 ;
	    RECT 139.1000 113.4000 140.2000 113.7000 ;
	    RECT 139.8000 111.1000 140.2000 113.4000 ;
	    RECT 140.6000 113.4000 141.7000 113.7000 ;
	    RECT 143.0000 113.4000 144.1000 113.7000 ;
	    RECT 145.4000 113.4000 146.5000 113.7000 ;
	    RECT 140.6000 111.1000 141.0000 113.4000 ;
	    RECT 143.0000 111.1000 143.4000 113.4000 ;
	    RECT 145.4000 111.1000 145.8000 113.4000 ;
	    RECT 2.2000 107.6000 2.6000 109.9000 ;
	    RECT 1.5000 107.3000 2.6000 107.6000 ;
	    RECT 3.0000 107.7000 3.4000 109.9000 ;
	    RECT 5.1000 109.2000 5.7000 109.9000 ;
	    RECT 5.1000 108.9000 5.8000 109.2000 ;
	    RECT 7.4000 108.9000 7.8000 109.9000 ;
	    RECT 9.6000 109.2000 10.0000 109.9000 ;
	    RECT 9.6000 108.9000 10.6000 109.2000 ;
	    RECT 5.4000 108.5000 5.8000 108.9000 ;
	    RECT 7.5000 108.6000 7.8000 108.9000 ;
	    RECT 7.5000 108.3000 8.9000 108.6000 ;
	    RECT 8.5000 108.2000 8.9000 108.3000 ;
	    RECT 9.4000 108.2000 9.8000 108.6000 ;
	    RECT 10.2000 108.5000 10.6000 108.9000 ;
	    RECT 6.2000 108.1000 6.6000 108.2000 ;
	    RECT 4.6000 107.8000 6.6000 108.1000 ;
	    RECT 4.5000 107.7000 5.0000 107.8000 ;
	    RECT 3.0000 107.4000 5.0000 107.7000 ;
	    RECT 1.5000 105.8000 1.8000 107.3000 ;
	    RECT 2.2000 106.1000 2.6000 106.6000 ;
	    RECT 3.0000 106.1000 3.4000 107.4000 ;
	    RECT 6.5000 107.1000 6.9000 107.2000 ;
	    RECT 9.4000 107.1000 9.7000 108.2000 ;
	    RECT 11.8000 107.5000 12.2000 109.9000 ;
	    RECT 12.6000 107.8000 13.0000 108.6000 ;
	    RECT 13.4000 108.1000 13.8000 109.9000 ;
	    RECT 15.0000 108.9000 15.4000 109.9000 ;
	    RECT 14.2000 108.1000 14.6000 108.6000 ;
	    RECT 13.4000 107.8000 14.6000 108.1000 ;
	    RECT 11.0000 107.1000 11.8000 107.2000 ;
	    RECT 6.3000 106.8000 11.8000 107.1000 ;
	    RECT 5.4000 106.4000 5.8000 106.5000 ;
	    RECT 2.2000 105.8000 3.4000 106.1000 ;
	    RECT 3.9000 106.1000 5.8000 106.4000 ;
	    RECT 6.3000 106.1000 6.6000 106.8000 ;
	    RECT 9.9000 106.7000 10.3000 106.8000 ;
	    RECT 9.4000 106.2000 9.8000 106.3000 ;
	    RECT 10.7000 106.2000 11.1000 106.3000 ;
	    RECT 7.0000 106.1000 7.4000 106.2000 ;
	    RECT 3.9000 106.0000 4.3000 106.1000 ;
	    RECT 6.2000 105.8000 7.4000 106.1000 ;
	    RECT 8.6000 105.9000 11.1000 106.2000 ;
	    RECT 8.6000 105.8000 9.0000 105.9000 ;
	    RECT 1.2000 105.4000 1.8000 105.8000 ;
	    RECT 1.5000 105.1000 1.8000 105.4000 ;
	    RECT 3.0000 105.7000 3.4000 105.8000 ;
	    RECT 4.7000 105.7000 5.1000 105.8000 ;
	    RECT 3.0000 105.4000 5.1000 105.7000 ;
	    RECT 1.5000 104.8000 2.6000 105.1000 ;
	    RECT 2.2000 101.1000 2.6000 104.8000 ;
	    RECT 3.0000 101.1000 3.4000 105.4000 ;
	    RECT 6.3000 105.2000 6.6000 105.8000 ;
	    RECT 9.4000 105.5000 12.2000 105.6000 ;
	    RECT 9.3000 105.4000 12.2000 105.5000 ;
	    RECT 5.4000 104.9000 6.6000 105.2000 ;
	    RECT 7.3000 105.3000 12.2000 105.4000 ;
	    RECT 7.3000 105.1000 9.7000 105.3000 ;
	    RECT 5.4000 104.4000 5.7000 104.9000 ;
	    RECT 5.0000 104.0000 5.7000 104.4000 ;
	    RECT 6.5000 104.5000 6.9000 104.6000 ;
	    RECT 7.3000 104.5000 7.6000 105.1000 ;
	    RECT 6.5000 104.2000 7.6000 104.5000 ;
	    RECT 7.9000 104.5000 10.6000 104.8000 ;
	    RECT 7.9000 104.4000 8.3000 104.5000 ;
	    RECT 10.2000 104.4000 10.6000 104.5000 ;
	    RECT 7.1000 103.7000 7.5000 103.8000 ;
	    RECT 8.5000 103.7000 8.9000 103.8000 ;
	    RECT 5.4000 103.1000 5.8000 103.5000 ;
	    RECT 7.1000 103.4000 8.9000 103.7000 ;
	    RECT 7.5000 103.1000 7.8000 103.4000 ;
	    RECT 10.2000 103.1000 10.6000 103.5000 ;
	    RECT 5.1000 101.1000 5.7000 103.1000 ;
	    RECT 7.4000 101.1000 7.8000 103.1000 ;
	    RECT 9.6000 102.8000 10.6000 103.1000 ;
	    RECT 9.6000 101.1000 10.0000 102.8000 ;
	    RECT 11.8000 101.1000 12.2000 105.3000 ;
	    RECT 13.4000 101.1000 13.8000 107.8000 ;
	    RECT 15.1000 107.2000 15.4000 108.9000 ;
	    RECT 18.2000 107.6000 18.6000 109.9000 ;
	    RECT 14.2000 106.8000 14.6000 107.2000 ;
	    RECT 15.0000 106.8000 15.4000 107.2000 ;
	    RECT 14.2000 106.1000 14.5000 106.8000 ;
	    RECT 15.1000 106.1000 15.4000 106.8000 ;
	    RECT 17.5000 107.3000 18.6000 107.6000 ;
	    RECT 19.0000 107.7000 19.4000 109.9000 ;
	    RECT 21.1000 109.2000 21.7000 109.9000 ;
	    RECT 21.1000 108.9000 21.8000 109.2000 ;
	    RECT 23.4000 108.9000 23.8000 109.9000 ;
	    RECT 25.6000 109.2000 26.0000 109.9000 ;
	    RECT 25.6000 108.9000 26.6000 109.2000 ;
	    RECT 21.4000 108.5000 21.8000 108.9000 ;
	    RECT 23.5000 108.6000 23.8000 108.9000 ;
	    RECT 23.5000 108.3000 24.9000 108.6000 ;
	    RECT 24.5000 108.2000 24.9000 108.3000 ;
	    RECT 25.4000 107.8000 25.8000 108.6000 ;
	    RECT 26.2000 108.5000 26.6000 108.9000 ;
	    RECT 20.5000 107.7000 20.9000 107.8000 ;
	    RECT 19.0000 107.4000 21.0000 107.7000 ;
	    RECT 14.2000 105.8000 15.4000 106.1000 ;
	    RECT 15.1000 105.1000 15.4000 105.8000 ;
	    RECT 15.8000 105.4000 16.2000 106.2000 ;
	    RECT 17.5000 105.8000 17.8000 107.3000 ;
	    RECT 18.2000 106.1000 18.6000 106.6000 ;
	    RECT 19.0000 106.1000 19.4000 107.4000 ;
	    RECT 20.6000 106.8000 21.0000 107.4000 ;
	    RECT 22.5000 107.1000 22.9000 107.2000 ;
	    RECT 25.4000 107.1000 25.7000 107.8000 ;
	    RECT 27.8000 107.5000 28.2000 109.9000 ;
	    RECT 28.6000 107.9000 29.0000 109.9000 ;
	    RECT 30.8000 108.1000 31.6000 109.9000 ;
	    RECT 28.6000 107.6000 29.8000 107.9000 ;
	    RECT 29.4000 107.5000 29.8000 107.6000 ;
	    RECT 30.1000 107.4000 30.5000 107.8000 ;
	    RECT 30.1000 107.2000 30.4000 107.4000 ;
	    RECT 27.0000 107.1000 27.8000 107.2000 ;
	    RECT 22.3000 106.8000 27.8000 107.1000 ;
	    RECT 28.6000 106.8000 29.4000 107.2000 ;
	    RECT 30.0000 106.8000 30.4000 107.2000 ;
	    RECT 21.4000 106.4000 21.8000 106.5000 ;
	    RECT 18.2000 105.8000 19.4000 106.1000 ;
	    RECT 19.9000 106.1000 21.8000 106.4000 ;
	    RECT 22.3000 106.1000 22.6000 106.8000 ;
	    RECT 25.9000 106.7000 26.3000 106.8000 ;
	    RECT 30.8000 106.4000 31.1000 108.1000 ;
	    RECT 33.4000 107.9000 33.8000 109.9000 ;
	    RECT 36.6000 108.9000 37.0000 109.9000 ;
	    RECT 38.2000 109.2000 38.6000 109.9000 ;
	    RECT 31.4000 107.7000 32.2000 107.8000 ;
	    RECT 31.4000 107.4000 32.4000 107.7000 ;
	    RECT 32.7000 107.6000 33.8000 107.9000 ;
	    RECT 36.4000 108.8000 37.0000 108.9000 ;
	    RECT 38.1000 108.8000 38.6000 109.2000 ;
	    RECT 36.4000 108.5000 38.4000 108.8000 ;
	    RECT 32.7000 107.5000 33.1000 107.6000 ;
	    RECT 32.1000 107.2000 32.4000 107.4000 ;
	    RECT 31.4000 106.7000 31.8000 107.1000 ;
	    RECT 32.1000 106.9000 33.8000 107.2000 ;
	    RECT 33.0000 106.8000 33.8000 106.9000 ;
	    RECT 25.4000 106.2000 25.8000 106.3000 ;
	    RECT 26.7000 106.2000 27.1000 106.3000 ;
	    RECT 30.6000 106.2000 31.1000 106.4000 ;
	    RECT 23.0000 106.1000 23.4000 106.2000 ;
	    RECT 19.9000 106.0000 20.3000 106.1000 ;
	    RECT 22.2000 105.8000 23.4000 106.1000 ;
	    RECT 24.6000 105.9000 27.1000 106.2000 ;
	    RECT 28.6000 106.1000 29.0000 106.2000 ;
	    RECT 30.2000 106.1000 31.1000 106.2000 ;
	    RECT 31.5000 106.4000 31.8000 106.7000 ;
	    RECT 31.5000 106.1000 32.8000 106.4000 ;
	    RECT 24.6000 105.8000 25.0000 105.9000 ;
	    RECT 28.6000 105.8000 30.9000 106.1000 ;
	    RECT 32.4000 106.0000 32.8000 106.1000 ;
	    RECT 17.2000 105.4000 17.8000 105.8000 ;
	    RECT 17.5000 105.1000 17.8000 105.4000 ;
	    RECT 19.0000 105.7000 19.4000 105.8000 ;
	    RECT 20.7000 105.7000 21.1000 105.8000 ;
	    RECT 19.0000 105.4000 21.1000 105.7000 ;
	    RECT 15.0000 104.7000 15.9000 105.1000 ;
	    RECT 17.5000 104.8000 18.6000 105.1000 ;
	    RECT 15.5000 101.1000 15.9000 104.7000 ;
	    RECT 18.2000 101.1000 18.6000 104.8000 ;
	    RECT 19.0000 101.1000 19.4000 105.4000 ;
	    RECT 22.3000 105.2000 22.6000 105.8000 ;
	    RECT 25.4000 105.5000 28.2000 105.6000 ;
	    RECT 25.3000 105.4000 28.2000 105.5000 ;
	    RECT 21.4000 104.9000 22.6000 105.2000 ;
	    RECT 23.3000 105.3000 28.2000 105.4000 ;
	    RECT 23.3000 105.1000 25.7000 105.3000 ;
	    RECT 21.4000 104.4000 21.7000 104.9000 ;
	    RECT 21.0000 104.0000 21.7000 104.4000 ;
	    RECT 22.5000 104.5000 22.9000 104.6000 ;
	    RECT 23.3000 104.5000 23.6000 105.1000 ;
	    RECT 22.5000 104.2000 23.6000 104.5000 ;
	    RECT 23.9000 104.5000 26.6000 104.8000 ;
	    RECT 23.9000 104.4000 24.3000 104.5000 ;
	    RECT 26.2000 104.4000 26.6000 104.5000 ;
	    RECT 23.1000 103.7000 23.5000 103.8000 ;
	    RECT 24.5000 103.7000 24.9000 103.8000 ;
	    RECT 21.4000 103.1000 21.8000 103.5000 ;
	    RECT 23.1000 103.4000 24.9000 103.7000 ;
	    RECT 23.5000 103.1000 23.8000 103.4000 ;
	    RECT 26.2000 103.1000 26.6000 103.5000 ;
	    RECT 21.1000 101.1000 21.7000 103.1000 ;
	    RECT 23.4000 101.1000 23.8000 103.1000 ;
	    RECT 25.6000 102.8000 26.6000 103.1000 ;
	    RECT 25.6000 101.1000 26.0000 102.8000 ;
	    RECT 27.8000 101.1000 28.2000 105.3000 ;
	    RECT 30.6000 105.1000 30.9000 105.8000 ;
	    RECT 31.3000 105.7000 31.7000 105.8000 ;
	    RECT 31.3000 105.4000 33.0000 105.7000 ;
	    RECT 32.7000 105.1000 33.0000 105.4000 ;
	    RECT 36.4000 105.2000 36.7000 108.5000 ;
	    RECT 38.5000 107.8000 39.4000 108.2000 ;
	    RECT 40.6000 107.8000 41.0000 108.6000 ;
	    RECT 37.8000 107.1000 38.6000 107.2000 ;
	    RECT 40.6000 107.1000 40.9000 107.8000 ;
	    RECT 37.8000 106.8000 40.9000 107.1000 ;
	    RECT 37.0000 106.1000 37.8000 106.2000 ;
	    RECT 40.6000 106.1000 41.0000 106.2000 ;
	    RECT 37.0000 105.8000 41.0000 106.1000 ;
	    RECT 28.6000 104.8000 29.8000 105.1000 ;
	    RECT 30.6000 104.8000 31.6000 105.1000 ;
	    RECT 28.6000 101.1000 29.0000 104.8000 ;
	    RECT 29.4000 104.7000 29.8000 104.8000 ;
	    RECT 30.8000 101.1000 31.6000 104.8000 ;
	    RECT 32.7000 104.8000 33.8000 105.1000 ;
	    RECT 35.0000 104.9000 36.7000 105.2000 ;
	    RECT 35.0000 104.8000 35.4000 104.9000 ;
	    RECT 32.7000 104.7000 33.1000 104.8000 ;
	    RECT 33.4000 101.1000 33.8000 104.8000 ;
	    RECT 35.1000 104.5000 35.4000 104.8000 ;
	    RECT 35.9000 104.5000 37.7000 104.6000 ;
	    RECT 34.2000 101.5000 34.6000 104.5000 ;
	    RECT 35.0000 101.7000 35.4000 104.5000 ;
	    RECT 35.8000 104.3000 37.7000 104.5000 ;
	    RECT 34.3000 101.4000 34.6000 101.5000 ;
	    RECT 35.8000 101.5000 36.2000 104.3000 ;
	    RECT 37.4000 104.1000 37.7000 104.3000 ;
	    RECT 38.3000 104.4000 40.1000 104.7000 ;
	    RECT 38.3000 104.1000 38.6000 104.4000 ;
	    RECT 35.8000 101.4000 36.1000 101.5000 ;
	    RECT 34.3000 101.1000 36.1000 101.4000 ;
	    RECT 36.6000 101.4000 37.0000 104.0000 ;
	    RECT 37.4000 101.7000 37.8000 104.1000 ;
	    RECT 38.2000 101.4000 38.6000 104.1000 ;
	    RECT 36.6000 101.1000 38.6000 101.4000 ;
	    RECT 39.8000 104.1000 40.1000 104.4000 ;
	    RECT 39.8000 101.1000 40.2000 104.1000 ;
	    RECT 41.4000 101.1000 41.8000 109.9000 ;
	    RECT 42.5000 109.2000 42.9000 109.9000 ;
	    RECT 42.2000 108.8000 42.9000 109.2000 ;
	    RECT 42.5000 108.4000 42.9000 108.8000 ;
	    RECT 42.2000 107.9000 42.9000 108.4000 ;
	    RECT 44.6000 107.9000 45.0000 109.9000 ;
	    RECT 45.4000 107.9000 45.8000 109.9000 ;
	    RECT 46.2000 108.0000 46.6000 109.9000 ;
	    RECT 47.8000 108.0000 48.2000 109.9000 ;
	    RECT 51.8000 109.2000 52.2000 109.9000 ;
	    RECT 51.8000 108.9000 52.3000 109.2000 ;
	    RECT 52.0000 108.8000 52.3000 108.9000 ;
	    RECT 53.4000 108.9000 53.8000 109.9000 ;
	    RECT 55.8000 109.1000 56.2000 109.2000 ;
	    RECT 56.6000 109.1000 57.0000 109.9000 ;
	    RECT 53.4000 108.8000 54.0000 108.9000 ;
	    RECT 55.8000 108.8000 57.0000 109.1000 ;
	    RECT 52.0000 108.5000 54.0000 108.8000 ;
	    RECT 46.2000 107.9000 48.2000 108.0000 ;
	    RECT 42.2000 106.2000 42.5000 107.9000 ;
	    RECT 44.6000 107.8000 44.9000 107.9000 ;
	    RECT 44.0000 107.6000 44.9000 107.8000 ;
	    RECT 42.8000 107.5000 44.9000 107.6000 ;
	    RECT 42.8000 107.3000 44.3000 107.5000 ;
	    RECT 42.8000 107.2000 43.2000 107.3000 ;
	    RECT 45.5000 107.2000 45.8000 107.9000 ;
	    RECT 46.3000 107.7000 48.1000 107.9000 ;
	    RECT 51.0000 107.8000 51.9000 108.2000 ;
	    RECT 47.4000 107.2000 47.8000 107.4000 ;
	    RECT 42.2000 105.8000 42.6000 106.2000 ;
	    RECT 42.2000 105.1000 42.5000 105.8000 ;
	    RECT 42.9000 105.5000 43.2000 107.2000 ;
	    RECT 44.6000 107.1000 45.0000 107.2000 ;
	    RECT 45.4000 107.1000 46.7000 107.2000 ;
	    RECT 43.6000 106.9000 44.0000 107.0000 ;
	    RECT 43.6000 106.6000 44.1000 106.9000 ;
	    RECT 43.8000 106.2000 44.1000 106.6000 ;
	    RECT 44.6000 106.8000 46.7000 107.1000 ;
	    RECT 47.4000 107.1000 48.2000 107.2000 ;
	    RECT 50.2000 107.1000 50.6000 107.2000 ;
	    RECT 47.4000 106.9000 50.6000 107.1000 ;
	    RECT 47.8000 106.8000 50.6000 106.9000 ;
	    RECT 51.8000 106.8000 52.6000 107.2000 ;
	    RECT 53.7000 107.1000 54.0000 108.5000 ;
	    RECT 56.6000 107.9000 57.0000 108.8000 ;
	    RECT 57.4000 108.0000 57.8000 109.9000 ;
	    RECT 59.0000 108.0000 59.4000 109.9000 ;
	    RECT 57.4000 107.9000 59.4000 108.0000 ;
	    RECT 59.8000 107.9000 60.2000 109.9000 ;
	    RECT 60.6000 108.0000 61.0000 109.9000 ;
	    RECT 62.2000 108.0000 62.6000 109.9000 ;
	    RECT 63.3000 109.2000 63.7000 109.9000 ;
	    RECT 63.0000 108.8000 63.7000 109.2000 ;
	    RECT 60.6000 107.9000 62.6000 108.0000 ;
	    RECT 63.3000 108.2000 63.7000 108.8000 ;
	    RECT 66.7000 108.2000 67.1000 109.9000 ;
	    RECT 63.3000 107.9000 64.2000 108.2000 ;
	    RECT 56.7000 107.2000 57.0000 107.9000 ;
	    RECT 57.5000 107.7000 59.3000 107.9000 ;
	    RECT 58.6000 107.2000 59.0000 107.4000 ;
	    RECT 59.9000 107.2000 60.2000 107.9000 ;
	    RECT 60.7000 107.7000 62.5000 107.9000 ;
	    RECT 61.8000 107.2000 62.2000 107.4000 ;
	    RECT 55.0000 107.1000 55.4000 107.2000 ;
	    RECT 53.7000 106.8000 55.4000 107.1000 ;
	    RECT 56.6000 106.8000 57.9000 107.2000 ;
	    RECT 58.6000 106.9000 59.4000 107.2000 ;
	    RECT 59.0000 106.8000 59.4000 106.9000 ;
	    RECT 59.8000 106.8000 61.1000 107.2000 ;
	    RECT 61.8000 106.9000 62.6000 107.2000 ;
	    RECT 62.2000 106.8000 62.6000 106.9000 ;
	    RECT 44.6000 106.4000 45.0000 106.8000 ;
	    RECT 43.8000 105.8000 44.2000 106.2000 ;
	    RECT 42.9000 105.2000 44.1000 105.5000 ;
	    RECT 42.2000 101.1000 42.6000 105.1000 ;
	    RECT 43.8000 103.1000 44.1000 105.2000 ;
	    RECT 45.4000 105.1000 45.8000 105.2000 ;
	    RECT 46.4000 105.1000 46.7000 106.8000 ;
	    RECT 47.0000 105.8000 47.4000 106.6000 ;
	    RECT 50.2000 106.1000 50.6000 106.2000 ;
	    RECT 52.6000 106.1000 53.4000 106.2000 ;
	    RECT 50.2000 105.8000 53.4000 106.1000 ;
	    RECT 53.7000 105.2000 54.0000 106.8000 ;
	    RECT 45.4000 104.8000 46.1000 105.1000 ;
	    RECT 46.4000 104.8000 46.9000 105.1000 ;
	    RECT 53.7000 104.9000 55.4000 105.2000 ;
	    RECT 45.8000 104.2000 46.1000 104.8000 ;
	    RECT 45.8000 103.8000 46.2000 104.2000 ;
	    RECT 43.8000 101.1000 44.2000 103.1000 ;
	    RECT 46.5000 101.1000 46.9000 104.8000 ;
	    RECT 55.0000 104.8000 55.4000 104.9000 ;
	    RECT 55.8000 105.1000 56.2000 105.2000 ;
	    RECT 56.6000 105.1000 57.0000 105.2000 ;
	    RECT 57.6000 105.1000 57.9000 106.8000 ;
	    RECT 58.2000 105.8000 58.6000 106.6000 ;
	    RECT 59.8000 105.1000 60.2000 105.2000 ;
	    RECT 60.8000 105.1000 61.1000 106.8000 ;
	    RECT 61.4000 106.1000 61.8000 106.6000 ;
	    RECT 62.2000 106.1000 62.6000 106.2000 ;
	    RECT 61.4000 105.8000 62.6000 106.1000 ;
	    RECT 55.8000 104.8000 57.3000 105.1000 ;
	    RECT 57.6000 104.8000 58.1000 105.1000 ;
	    RECT 59.8000 104.8000 60.5000 105.1000 ;
	    RECT 60.8000 104.8000 61.3000 105.1000 ;
	    RECT 50.3000 104.4000 52.1000 104.7000 ;
	    RECT 50.3000 104.1000 50.6000 104.4000 ;
	    RECT 50.2000 101.1000 50.6000 104.1000 ;
	    RECT 51.8000 104.1000 52.1000 104.4000 ;
	    RECT 52.7000 104.5000 54.5000 104.6000 ;
	    RECT 55.0000 104.5000 55.3000 104.8000 ;
	    RECT 52.7000 104.3000 54.6000 104.5000 ;
	    RECT 52.7000 104.1000 53.0000 104.3000 ;
	    RECT 51.8000 101.4000 52.2000 104.1000 ;
	    RECT 52.6000 101.7000 53.0000 104.1000 ;
	    RECT 53.4000 101.4000 53.8000 104.0000 ;
	    RECT 54.2000 101.5000 54.6000 104.3000 ;
	    RECT 55.0000 101.7000 55.4000 104.5000 ;
	    RECT 51.8000 101.1000 53.8000 101.4000 ;
	    RECT 54.3000 101.4000 54.6000 101.5000 ;
	    RECT 55.8000 101.5000 56.2000 104.5000 ;
	    RECT 57.0000 104.2000 57.3000 104.8000 ;
	    RECT 57.0000 103.8000 57.4000 104.2000 ;
	    RECT 55.8000 101.4000 56.1000 101.5000 ;
	    RECT 54.3000 101.1000 56.1000 101.4000 ;
	    RECT 57.7000 101.1000 58.1000 104.8000 ;
	    RECT 60.2000 104.2000 60.5000 104.8000 ;
	    RECT 60.2000 103.8000 60.6000 104.2000 ;
	    RECT 60.9000 101.1000 61.3000 104.8000 ;
	    RECT 63.0000 104.4000 63.4000 105.2000 ;
	    RECT 63.8000 101.1000 64.2000 107.9000 ;
	    RECT 66.2000 107.9000 67.1000 108.2000 ;
	    RECT 67.8000 107.9000 68.2000 109.9000 ;
	    RECT 70.0000 108.1000 70.8000 109.9000 ;
	    RECT 64.6000 106.8000 65.0000 107.6000 ;
	    RECT 65.4000 106.8000 65.8000 107.6000 ;
	    RECT 64.6000 106.1000 64.9000 106.8000 ;
	    RECT 66.2000 106.1000 66.6000 107.9000 ;
	    RECT 67.8000 107.6000 68.9000 107.9000 ;
	    RECT 69.4000 107.7000 70.2000 107.8000 ;
	    RECT 68.5000 107.5000 68.9000 107.6000 ;
	    RECT 69.2000 107.4000 70.2000 107.7000 ;
	    RECT 69.2000 107.2000 69.5000 107.4000 ;
	    RECT 67.0000 107.1000 67.4000 107.2000 ;
	    RECT 67.8000 107.1000 69.5000 107.2000 ;
	    RECT 67.0000 106.9000 69.5000 107.1000 ;
	    RECT 67.0000 106.8000 68.6000 106.9000 ;
	    RECT 69.8000 106.7000 70.2000 107.1000 ;
	    RECT 69.8000 106.4000 70.1000 106.7000 ;
	    RECT 64.6000 105.8000 66.6000 106.1000 ;
	    RECT 68.8000 106.1000 70.1000 106.4000 ;
	    RECT 70.5000 106.4000 70.8000 108.1000 ;
	    RECT 72.6000 107.9000 73.0000 109.9000 ;
	    RECT 71.1000 107.4000 71.5000 107.8000 ;
	    RECT 71.8000 107.6000 73.0000 107.9000 ;
	    RECT 71.8000 107.5000 72.2000 107.6000 ;
	    RECT 71.2000 107.2000 71.5000 107.4000 ;
	    RECT 71.2000 106.8000 71.6000 107.2000 ;
	    RECT 72.2000 107.1000 73.0000 107.2000 ;
	    RECT 73.4000 107.1000 73.8000 109.9000 ;
	    RECT 74.2000 107.8000 74.6000 108.6000 ;
	    RECT 72.2000 106.8000 73.8000 107.1000 ;
	    RECT 70.5000 106.2000 71.0000 106.4000 ;
	    RECT 70.5000 106.1000 71.4000 106.2000 ;
	    RECT 72.6000 106.1000 73.0000 106.2000 ;
	    RECT 68.8000 106.0000 69.2000 106.1000 ;
	    RECT 70.7000 105.8000 73.0000 106.1000 ;
	    RECT 65.4000 104.1000 65.8000 104.2000 ;
	    RECT 66.2000 104.1000 66.6000 105.8000 ;
	    RECT 69.9000 105.7000 70.3000 105.8000 ;
	    RECT 68.6000 105.4000 70.3000 105.7000 ;
	    RECT 67.0000 104.4000 67.4000 105.2000 ;
	    RECT 68.6000 105.1000 68.9000 105.4000 ;
	    RECT 70.7000 105.1000 71.0000 105.8000 ;
	    RECT 67.8000 104.8000 68.9000 105.1000 ;
	    RECT 65.4000 103.8000 66.6000 104.1000 ;
	    RECT 66.2000 101.1000 66.6000 103.8000 ;
	    RECT 67.8000 101.1000 68.2000 104.8000 ;
	    RECT 68.5000 104.7000 68.9000 104.8000 ;
	    RECT 70.0000 104.8000 71.0000 105.1000 ;
	    RECT 71.8000 104.8000 73.0000 105.1000 ;
	    RECT 70.0000 101.1000 70.8000 104.8000 ;
	    RECT 71.8000 104.7000 72.2000 104.8000 ;
	    RECT 72.6000 101.1000 73.0000 104.8000 ;
	    RECT 73.4000 101.1000 73.8000 106.8000 ;
	    RECT 75.0000 107.7000 75.4000 109.9000 ;
	    RECT 77.1000 109.2000 77.7000 109.9000 ;
	    RECT 77.1000 108.9000 77.8000 109.2000 ;
	    RECT 79.4000 108.9000 79.8000 109.9000 ;
	    RECT 81.6000 109.2000 82.0000 109.9000 ;
	    RECT 81.6000 108.9000 82.6000 109.2000 ;
	    RECT 77.4000 108.5000 77.8000 108.9000 ;
	    RECT 79.5000 108.6000 79.8000 108.9000 ;
	    RECT 79.5000 108.3000 80.9000 108.6000 ;
	    RECT 80.5000 108.2000 80.9000 108.3000 ;
	    RECT 81.4000 108.2000 81.8000 108.6000 ;
	    RECT 82.2000 108.5000 82.6000 108.9000 ;
	    RECT 76.5000 107.7000 76.9000 107.8000 ;
	    RECT 75.0000 107.4000 76.9000 107.7000 ;
	    RECT 75.0000 105.7000 75.4000 107.4000 ;
	    RECT 78.5000 107.1000 78.9000 107.2000 ;
	    RECT 81.4000 107.1000 81.7000 108.2000 ;
	    RECT 83.8000 107.5000 84.2000 109.9000 ;
	    RECT 84.6000 107.6000 85.0000 109.9000 ;
	    RECT 84.6000 107.3000 85.7000 107.6000 ;
	    RECT 87.0000 107.5000 87.4000 109.9000 ;
	    RECT 89.2000 109.2000 89.6000 109.9000 ;
	    RECT 88.6000 108.9000 89.6000 109.2000 ;
	    RECT 91.4000 108.9000 91.8000 109.9000 ;
	    RECT 93.5000 109.2000 94.1000 109.9000 ;
	    RECT 93.4000 108.9000 94.1000 109.2000 ;
	    RECT 88.6000 108.5000 89.0000 108.9000 ;
	    RECT 91.4000 108.6000 91.7000 108.9000 ;
	    RECT 89.4000 108.2000 89.8000 108.6000 ;
	    RECT 90.3000 108.3000 91.7000 108.6000 ;
	    RECT 93.4000 108.5000 93.8000 108.9000 ;
	    RECT 90.3000 108.2000 90.7000 108.3000 ;
	    RECT 83.0000 107.1000 83.8000 107.2000 ;
	    RECT 78.3000 106.8000 83.8000 107.1000 ;
	    RECT 77.4000 106.4000 77.8000 106.5000 ;
	    RECT 75.9000 106.1000 77.8000 106.4000 ;
	    RECT 78.3000 106.2000 78.6000 106.8000 ;
	    RECT 81.9000 106.7000 82.3000 106.8000 ;
	    RECT 82.7000 106.2000 83.1000 106.3000 ;
	    RECT 75.9000 106.0000 76.3000 106.1000 ;
	    RECT 78.2000 105.8000 78.6000 106.2000 ;
	    RECT 80.6000 105.9000 83.1000 106.2000 ;
	    RECT 80.6000 105.8000 81.0000 105.9000 ;
	    RECT 84.6000 105.8000 85.0000 106.6000 ;
	    RECT 85.4000 105.8000 85.7000 107.3000 ;
	    RECT 87.4000 107.1000 88.2000 107.2000 ;
	    RECT 89.5000 107.1000 89.8000 108.2000 ;
	    RECT 92.6000 107.8000 93.0000 108.2000 ;
	    RECT 92.6000 107.2000 92.9000 107.8000 ;
	    RECT 94.3000 107.7000 94.7000 107.8000 ;
	    RECT 95.8000 107.7000 96.2000 109.9000 ;
	    RECT 94.3000 107.4000 96.2000 107.7000 ;
	    RECT 98.2000 107.5000 98.6000 109.9000 ;
	    RECT 100.4000 109.2000 100.8000 109.9000 ;
	    RECT 99.8000 108.9000 100.8000 109.2000 ;
	    RECT 102.6000 108.9000 103.0000 109.9000 ;
	    RECT 104.7000 109.2000 105.3000 109.9000 ;
	    RECT 104.6000 108.9000 105.3000 109.2000 ;
	    RECT 99.8000 108.5000 100.2000 108.9000 ;
	    RECT 102.6000 108.6000 102.9000 108.9000 ;
	    RECT 100.6000 108.2000 101.0000 108.6000 ;
	    RECT 101.5000 108.3000 102.9000 108.6000 ;
	    RECT 104.6000 108.5000 105.0000 108.9000 ;
	    RECT 101.5000 108.2000 101.9000 108.3000 ;
	    RECT 92.3000 107.1000 92.9000 107.2000 ;
	    RECT 87.4000 106.8000 92.9000 107.1000 ;
	    RECT 88.9000 106.7000 89.3000 106.8000 ;
	    RECT 88.1000 106.2000 88.5000 106.3000 ;
	    RECT 89.4000 106.2000 89.8000 106.3000 ;
	    RECT 88.1000 105.9000 90.6000 106.2000 ;
	    RECT 90.2000 105.8000 90.6000 105.9000 ;
	    RECT 76.7000 105.7000 77.1000 105.8000 ;
	    RECT 75.0000 105.4000 77.1000 105.7000 ;
	    RECT 74.2000 104.1000 74.6000 104.2000 ;
	    RECT 75.0000 104.1000 75.4000 105.4000 ;
	    RECT 78.3000 105.2000 78.6000 105.8000 ;
	    RECT 81.4000 105.5000 84.2000 105.6000 ;
	    RECT 81.3000 105.4000 84.2000 105.5000 ;
	    RECT 77.4000 104.9000 78.6000 105.2000 ;
	    RECT 79.3000 105.3000 84.2000 105.4000 ;
	    RECT 79.3000 105.1000 81.7000 105.3000 ;
	    RECT 77.4000 104.4000 77.7000 104.9000 ;
	    RECT 74.2000 103.8000 75.4000 104.1000 ;
	    RECT 77.0000 104.0000 77.7000 104.4000 ;
	    RECT 78.5000 104.5000 78.9000 104.6000 ;
	    RECT 79.3000 104.5000 79.6000 105.1000 ;
	    RECT 78.5000 104.2000 79.6000 104.5000 ;
	    RECT 79.9000 104.5000 82.6000 104.8000 ;
	    RECT 79.9000 104.4000 80.3000 104.5000 ;
	    RECT 82.2000 104.4000 82.6000 104.5000 ;
	    RECT 75.0000 101.1000 75.4000 103.8000 ;
	    RECT 79.1000 103.7000 79.5000 103.8000 ;
	    RECT 80.5000 103.7000 80.9000 103.8000 ;
	    RECT 77.4000 103.1000 77.8000 103.5000 ;
	    RECT 79.1000 103.4000 80.9000 103.7000 ;
	    RECT 79.5000 103.1000 79.8000 103.4000 ;
	    RECT 82.2000 103.1000 82.6000 103.5000 ;
	    RECT 77.1000 101.1000 77.7000 103.1000 ;
	    RECT 79.4000 101.1000 79.8000 103.1000 ;
	    RECT 81.6000 102.8000 82.6000 103.1000 ;
	    RECT 81.6000 101.1000 82.0000 102.8000 ;
	    RECT 83.8000 101.1000 84.2000 105.3000 ;
	    RECT 85.4000 105.4000 86.0000 105.8000 ;
	    RECT 87.0000 105.5000 89.8000 105.6000 ;
	    RECT 87.0000 105.4000 89.9000 105.5000 ;
	    RECT 85.4000 105.1000 85.7000 105.4000 ;
	    RECT 84.6000 104.8000 85.7000 105.1000 ;
	    RECT 87.0000 105.3000 91.9000 105.4000 ;
	    RECT 84.6000 101.1000 85.0000 104.8000 ;
	    RECT 87.0000 101.1000 87.4000 105.3000 ;
	    RECT 89.5000 105.1000 91.9000 105.3000 ;
	    RECT 88.6000 104.5000 91.3000 104.8000 ;
	    RECT 88.6000 104.4000 89.0000 104.5000 ;
	    RECT 90.9000 104.4000 91.3000 104.5000 ;
	    RECT 91.6000 104.5000 91.9000 105.1000 ;
	    RECT 92.6000 105.2000 92.9000 106.8000 ;
	    RECT 93.4000 106.4000 93.8000 106.5000 ;
	    RECT 93.4000 106.1000 95.3000 106.4000 ;
	    RECT 94.9000 106.0000 95.3000 106.1000 ;
	    RECT 94.1000 105.7000 94.5000 105.8000 ;
	    RECT 95.8000 105.7000 96.2000 107.4000 ;
	    RECT 98.6000 107.1000 99.4000 107.2000 ;
	    RECT 100.7000 107.1000 101.0000 108.2000 ;
	    RECT 105.5000 107.7000 105.9000 107.8000 ;
	    RECT 107.0000 107.7000 107.4000 109.9000 ;
	    RECT 107.8000 107.8000 108.2000 108.6000 ;
	    RECT 105.5000 107.4000 107.4000 107.7000 ;
	    RECT 103.5000 107.1000 103.9000 107.2000 ;
	    RECT 98.6000 106.8000 104.1000 107.1000 ;
	    RECT 100.1000 106.7000 100.5000 106.8000 ;
	    RECT 99.3000 106.2000 99.7000 106.3000 ;
	    RECT 99.3000 105.9000 101.8000 106.2000 ;
	    RECT 101.4000 105.8000 101.8000 105.9000 ;
	    RECT 94.1000 105.4000 96.2000 105.7000 ;
	    RECT 92.6000 104.9000 93.8000 105.2000 ;
	    RECT 92.3000 104.5000 92.7000 104.6000 ;
	    RECT 91.6000 104.2000 92.7000 104.5000 ;
	    RECT 93.5000 104.4000 93.8000 104.9000 ;
	    RECT 93.5000 104.0000 94.2000 104.4000 ;
	    RECT 90.3000 103.7000 90.7000 103.8000 ;
	    RECT 91.7000 103.7000 92.1000 103.8000 ;
	    RECT 88.6000 103.1000 89.0000 103.5000 ;
	    RECT 90.3000 103.4000 92.1000 103.7000 ;
	    RECT 91.4000 103.1000 91.7000 103.4000 ;
	    RECT 93.4000 103.1000 93.8000 103.5000 ;
	    RECT 88.6000 102.8000 89.6000 103.1000 ;
	    RECT 89.2000 101.1000 89.6000 102.8000 ;
	    RECT 91.4000 101.1000 91.8000 103.1000 ;
	    RECT 93.5000 101.1000 94.1000 103.1000 ;
	    RECT 95.8000 101.1000 96.2000 105.4000 ;
	    RECT 98.2000 105.5000 101.0000 105.6000 ;
	    RECT 98.2000 105.4000 101.1000 105.5000 ;
	    RECT 98.2000 105.3000 103.1000 105.4000 ;
	    RECT 98.2000 101.1000 98.6000 105.3000 ;
	    RECT 100.7000 105.1000 103.1000 105.3000 ;
	    RECT 99.8000 104.5000 102.5000 104.8000 ;
	    RECT 99.8000 104.4000 100.2000 104.5000 ;
	    RECT 102.1000 104.4000 102.5000 104.5000 ;
	    RECT 102.8000 104.5000 103.1000 105.1000 ;
	    RECT 103.8000 105.2000 104.1000 106.8000 ;
	    RECT 104.6000 106.4000 105.0000 106.5000 ;
	    RECT 104.6000 106.1000 106.5000 106.4000 ;
	    RECT 106.1000 106.0000 106.5000 106.1000 ;
	    RECT 105.3000 105.7000 105.7000 105.8000 ;
	    RECT 107.0000 105.7000 107.4000 107.4000 ;
	    RECT 105.3000 105.4000 107.4000 105.7000 ;
	    RECT 103.8000 104.9000 105.0000 105.2000 ;
	    RECT 103.5000 104.5000 103.9000 104.6000 ;
	    RECT 102.8000 104.2000 103.9000 104.5000 ;
	    RECT 104.7000 104.4000 105.0000 104.9000 ;
	    RECT 104.7000 104.0000 105.4000 104.4000 ;
	    RECT 101.5000 103.7000 101.9000 103.8000 ;
	    RECT 102.9000 103.7000 103.3000 103.8000 ;
	    RECT 99.8000 103.1000 100.2000 103.5000 ;
	    RECT 101.5000 103.4000 103.3000 103.7000 ;
	    RECT 102.6000 103.1000 102.9000 103.4000 ;
	    RECT 104.6000 103.1000 105.0000 103.5000 ;
	    RECT 99.8000 102.8000 100.8000 103.1000 ;
	    RECT 100.4000 101.1000 100.8000 102.8000 ;
	    RECT 102.6000 101.1000 103.0000 103.1000 ;
	    RECT 104.7000 101.1000 105.3000 103.1000 ;
	    RECT 107.0000 101.1000 107.4000 105.4000 ;
	    RECT 108.6000 101.1000 109.0000 109.9000 ;
	    RECT 109.4000 108.5000 109.8000 109.5000 ;
	    RECT 109.4000 107.4000 109.7000 108.5000 ;
	    RECT 111.5000 108.0000 111.9000 109.5000 ;
	    RECT 111.5000 107.7000 112.3000 108.0000 ;
	    RECT 114.2000 107.9000 114.6000 109.9000 ;
	    RECT 115.0000 108.0000 115.4000 109.9000 ;
	    RECT 116.6000 108.0000 117.0000 109.9000 ;
	    RECT 115.0000 107.9000 117.0000 108.0000 ;
	    RECT 117.4000 108.5000 117.8000 109.5000 ;
	    RECT 111.9000 107.5000 112.3000 107.7000 ;
	    RECT 109.4000 107.1000 111.5000 107.4000 ;
	    RECT 111.0000 106.9000 111.5000 107.1000 ;
	    RECT 112.0000 107.2000 112.3000 107.5000 ;
	    RECT 114.3000 107.2000 114.6000 107.9000 ;
	    RECT 115.1000 107.7000 116.9000 107.9000 ;
	    RECT 117.4000 107.4000 117.7000 108.5000 ;
	    RECT 119.5000 108.0000 119.9000 109.5000 ;
	    RECT 119.5000 107.7000 120.3000 108.0000 ;
	    RECT 119.9000 107.5000 120.3000 107.7000 ;
	    RECT 116.2000 107.2000 116.6000 107.4000 ;
	    RECT 109.4000 105.8000 109.8000 106.6000 ;
	    RECT 111.0000 106.5000 111.7000 106.9000 ;
	    RECT 112.0000 106.8000 113.0000 107.2000 ;
	    RECT 114.2000 106.8000 115.5000 107.2000 ;
	    RECT 116.2000 106.9000 117.0000 107.2000 ;
	    RECT 117.4000 107.1000 119.5000 107.4000 ;
	    RECT 116.6000 106.8000 117.0000 106.9000 ;
	    RECT 119.0000 106.9000 119.5000 107.1000 ;
	    RECT 120.0000 107.2000 120.3000 107.5000 ;
	    RECT 123.8000 107.9000 124.2000 109.9000 ;
	    RECT 126.2000 108.9000 126.6000 109.9000 ;
	    RECT 124.5000 108.2000 124.9000 108.6000 ;
	    RECT 111.0000 105.5000 111.3000 106.5000 ;
	    RECT 109.4000 105.2000 111.3000 105.5000 ;
	    RECT 109.4000 103.5000 109.7000 105.2000 ;
	    RECT 112.0000 104.9000 112.3000 106.8000 ;
	    RECT 112.6000 106.1000 113.0000 106.2000 ;
	    RECT 115.2000 106.1000 115.5000 106.8000 ;
	    RECT 112.6000 105.8000 115.5000 106.1000 ;
	    RECT 115.8000 105.8000 116.2000 106.6000 ;
	    RECT 117.4000 105.8000 117.8000 106.6000 ;
	    RECT 119.0000 106.5000 119.7000 106.9000 ;
	    RECT 120.0000 106.8000 121.0000 107.2000 ;
	    RECT 121.4000 107.1000 121.8000 107.2000 ;
	    RECT 123.0000 107.1000 123.4000 107.2000 ;
	    RECT 121.4000 106.8000 123.4000 107.1000 ;
	    RECT 112.6000 105.4000 113.0000 105.8000 ;
	    RECT 111.5000 104.6000 112.3000 104.9000 ;
	    RECT 114.2000 105.1000 114.6000 105.2000 ;
	    RECT 115.2000 105.1000 115.5000 105.8000 ;
	    RECT 119.0000 105.5000 119.3000 106.5000 ;
	    RECT 117.4000 105.2000 119.3000 105.5000 ;
	    RECT 114.2000 104.8000 114.9000 105.1000 ;
	    RECT 115.2000 104.8000 115.7000 105.1000 ;
	    RECT 109.4000 101.5000 109.8000 103.5000 ;
	    RECT 111.5000 102.2000 111.9000 104.6000 ;
	    RECT 114.6000 104.2000 114.9000 104.8000 ;
	    RECT 114.6000 103.8000 115.0000 104.2000 ;
	    RECT 111.0000 101.8000 111.9000 102.2000 ;
	    RECT 111.5000 101.1000 111.9000 101.8000 ;
	    RECT 115.3000 101.1000 115.7000 104.8000 ;
	    RECT 117.4000 103.5000 117.7000 105.2000 ;
	    RECT 120.0000 104.9000 120.3000 106.8000 ;
	    RECT 123.0000 106.4000 123.4000 106.8000 ;
	    RECT 120.6000 105.4000 121.0000 106.2000 ;
	    RECT 122.2000 106.1000 122.6000 106.2000 ;
	    RECT 123.8000 106.1000 124.1000 107.9000 ;
	    RECT 124.6000 107.8000 125.0000 108.2000 ;
	    RECT 125.4000 107.8000 125.8000 108.6000 ;
	    RECT 124.6000 107.1000 124.9000 107.8000 ;
	    RECT 126.3000 107.2000 126.6000 108.9000 ;
	    RECT 127.8000 108.0000 128.2000 109.9000 ;
	    RECT 129.4000 108.0000 129.8000 109.9000 ;
	    RECT 127.8000 107.9000 129.8000 108.0000 ;
	    RECT 130.2000 107.9000 130.6000 109.9000 ;
	    RECT 132.6000 107.9000 133.0000 109.9000 ;
	    RECT 135.0000 108.9000 135.4000 109.9000 ;
	    RECT 133.3000 108.2000 133.7000 108.6000 ;
	    RECT 127.9000 107.7000 129.7000 107.9000 ;
	    RECT 128.2000 107.2000 128.6000 107.4000 ;
	    RECT 130.2000 107.2000 130.5000 107.9000 ;
	    RECT 126.2000 107.1000 126.6000 107.2000 ;
	    RECT 124.6000 106.8000 126.6000 107.1000 ;
	    RECT 127.8000 106.9000 128.6000 107.2000 ;
	    RECT 127.8000 106.8000 128.2000 106.9000 ;
	    RECT 129.3000 106.8000 130.6000 107.2000 ;
	    RECT 124.6000 106.1000 125.0000 106.2000 ;
	    RECT 122.2000 105.8000 123.0000 106.1000 ;
	    RECT 123.8000 105.8000 125.0000 106.1000 ;
	    RECT 122.6000 105.6000 123.0000 105.8000 ;
	    RECT 124.6000 105.1000 124.9000 105.8000 ;
	    RECT 126.3000 105.1000 126.6000 106.8000 ;
	    RECT 127.0000 105.4000 127.4000 106.2000 ;
	    RECT 128.6000 105.8000 129.0000 106.6000 ;
	    RECT 129.3000 105.1000 129.6000 106.8000 ;
	    RECT 131.8000 106.4000 132.2000 107.2000 ;
	    RECT 131.0000 106.1000 131.4000 106.2000 ;
	    RECT 132.6000 106.1000 132.9000 107.9000 ;
	    RECT 133.4000 107.8000 133.8000 108.2000 ;
	    RECT 134.2000 107.8000 134.6000 108.6000 ;
	    RECT 133.4000 107.1000 133.7000 107.8000 ;
	    RECT 135.1000 107.2000 135.4000 108.9000 ;
	    RECT 135.0000 107.1000 135.4000 107.2000 ;
	    RECT 133.4000 106.8000 135.4000 107.1000 ;
	    RECT 133.4000 106.1000 133.8000 106.2000 ;
	    RECT 131.0000 105.8000 131.8000 106.1000 ;
	    RECT 132.6000 105.8000 133.8000 106.1000 ;
	    RECT 131.4000 105.6000 131.8000 105.8000 ;
	    RECT 130.2000 105.1000 130.6000 105.2000 ;
	    RECT 133.4000 105.1000 133.7000 105.8000 ;
	    RECT 135.1000 105.1000 135.4000 106.8000 ;
	    RECT 137.4000 108.9000 137.8000 109.9000 ;
	    RECT 137.4000 107.2000 137.7000 108.9000 ;
	    RECT 138.2000 107.8000 138.6000 108.6000 ;
	    RECT 139.0000 107.5000 139.4000 109.9000 ;
	    RECT 141.2000 109.2000 141.6000 109.9000 ;
	    RECT 140.6000 108.9000 141.6000 109.2000 ;
	    RECT 143.4000 108.9000 143.8000 109.9000 ;
	    RECT 145.5000 109.2000 146.1000 109.9000 ;
	    RECT 145.4000 108.9000 146.1000 109.2000 ;
	    RECT 140.6000 108.5000 141.0000 108.9000 ;
	    RECT 143.4000 108.6000 143.7000 108.9000 ;
	    RECT 141.4000 108.2000 141.8000 108.6000 ;
	    RECT 142.3000 108.3000 143.7000 108.6000 ;
	    RECT 145.4000 108.5000 145.8000 108.9000 ;
	    RECT 142.3000 108.2000 142.7000 108.3000 ;
	    RECT 137.4000 106.8000 137.8000 107.2000 ;
	    RECT 139.4000 107.1000 140.2000 107.2000 ;
	    RECT 141.5000 107.1000 141.8000 108.2000 ;
	    RECT 146.3000 107.7000 146.7000 107.8000 ;
	    RECT 147.8000 107.7000 148.2000 109.9000 ;
	    RECT 146.3000 107.4000 148.2000 107.7000 ;
	    RECT 144.3000 107.1000 144.7000 107.2000 ;
	    RECT 139.4000 106.8000 144.9000 107.1000 ;
	    RECT 135.8000 106.1000 136.2000 106.2000 ;
	    RECT 136.6000 106.1000 137.0000 106.2000 ;
	    RECT 135.8000 105.8000 137.0000 106.1000 ;
	    RECT 135.8000 105.4000 136.2000 105.8000 ;
	    RECT 136.6000 105.4000 137.0000 105.8000 ;
	    RECT 137.4000 106.1000 137.7000 106.8000 ;
	    RECT 140.9000 106.7000 141.3000 106.8000 ;
	    RECT 140.1000 106.2000 140.5000 106.3000 ;
	    RECT 138.2000 106.1000 138.6000 106.2000 ;
	    RECT 137.4000 105.8000 138.6000 106.1000 ;
	    RECT 140.1000 105.9000 142.6000 106.2000 ;
	    RECT 142.2000 105.8000 142.6000 105.9000 ;
	    RECT 137.4000 105.1000 137.7000 105.8000 ;
	    RECT 139.0000 105.5000 141.8000 105.6000 ;
	    RECT 139.0000 105.4000 141.9000 105.5000 ;
	    RECT 139.0000 105.3000 143.9000 105.4000 ;
	    RECT 119.5000 104.6000 120.3000 104.9000 ;
	    RECT 122.2000 104.8000 124.2000 105.1000 ;
	    RECT 117.4000 101.5000 117.8000 103.5000 ;
	    RECT 119.5000 102.2000 119.9000 104.6000 ;
	    RECT 119.0000 101.8000 119.9000 102.2000 ;
	    RECT 119.5000 101.1000 119.9000 101.8000 ;
	    RECT 122.2000 101.1000 122.6000 104.8000 ;
	    RECT 123.8000 101.1000 124.2000 104.8000 ;
	    RECT 124.6000 101.1000 125.0000 105.1000 ;
	    RECT 126.2000 104.7000 127.1000 105.1000 ;
	    RECT 126.7000 101.1000 127.1000 104.7000 ;
	    RECT 129.1000 104.8000 129.6000 105.1000 ;
	    RECT 129.9000 104.8000 130.6000 105.1000 ;
	    RECT 131.0000 104.8000 133.0000 105.1000 ;
	    RECT 129.1000 104.2000 129.5000 104.8000 ;
	    RECT 129.9000 104.2000 130.2000 104.8000 ;
	    RECT 128.6000 103.8000 129.5000 104.2000 ;
	    RECT 129.8000 103.8000 130.2000 104.2000 ;
	    RECT 129.1000 101.1000 129.5000 103.8000 ;
	    RECT 131.0000 101.1000 131.4000 104.8000 ;
	    RECT 132.6000 101.1000 133.0000 104.8000 ;
	    RECT 133.4000 101.1000 133.8000 105.1000 ;
	    RECT 135.0000 104.7000 135.9000 105.1000 ;
	    RECT 135.5000 101.1000 135.9000 104.7000 ;
	    RECT 136.9000 104.7000 137.8000 105.1000 ;
	    RECT 136.9000 101.1000 137.3000 104.7000 ;
	    RECT 139.0000 101.1000 139.4000 105.3000 ;
	    RECT 141.5000 105.1000 143.9000 105.3000 ;
	    RECT 140.6000 104.5000 143.3000 104.8000 ;
	    RECT 140.6000 104.4000 141.0000 104.5000 ;
	    RECT 142.9000 104.4000 143.3000 104.5000 ;
	    RECT 143.6000 104.5000 143.9000 105.1000 ;
	    RECT 144.6000 105.2000 144.9000 106.8000 ;
	    RECT 145.4000 106.4000 145.8000 106.5000 ;
	    RECT 145.4000 106.1000 147.3000 106.4000 ;
	    RECT 146.9000 106.0000 147.3000 106.1000 ;
	    RECT 146.1000 105.7000 146.5000 105.8000 ;
	    RECT 147.8000 105.7000 148.2000 107.4000 ;
	    RECT 146.1000 105.4000 148.2000 105.7000 ;
	    RECT 144.6000 104.9000 145.8000 105.2000 ;
	    RECT 144.3000 104.5000 144.7000 104.6000 ;
	    RECT 143.6000 104.2000 144.7000 104.5000 ;
	    RECT 145.5000 104.4000 145.8000 104.9000 ;
	    RECT 145.5000 104.0000 146.2000 104.4000 ;
	    RECT 142.3000 103.7000 142.7000 103.8000 ;
	    RECT 143.7000 103.7000 144.1000 103.8000 ;
	    RECT 140.6000 103.1000 141.0000 103.5000 ;
	    RECT 142.3000 103.4000 144.1000 103.7000 ;
	    RECT 143.4000 103.1000 143.7000 103.4000 ;
	    RECT 145.4000 103.1000 145.8000 103.5000 ;
	    RECT 140.6000 102.8000 141.6000 103.1000 ;
	    RECT 141.2000 101.1000 141.6000 102.8000 ;
	    RECT 143.4000 101.1000 143.8000 103.1000 ;
	    RECT 145.5000 101.1000 146.1000 103.1000 ;
	    RECT 147.8000 101.1000 148.2000 105.4000 ;
	    RECT 2.2000 96.2000 2.6000 99.9000 ;
	    RECT 4.6000 96.2000 5.0000 99.9000 ;
	    RECT 1.5000 95.9000 2.6000 96.2000 ;
	    RECT 3.9000 95.9000 5.0000 96.2000 ;
	    RECT 1.5000 95.6000 1.8000 95.9000 ;
	    RECT 3.9000 95.6000 4.2000 95.9000 ;
	    RECT 1.2000 95.2000 1.8000 95.6000 ;
	    RECT 3.6000 95.2000 4.2000 95.6000 ;
	    RECT 5.4000 95.6000 5.8000 99.9000 ;
	    RECT 7.5000 97.9000 8.1000 99.9000 ;
	    RECT 9.8000 97.9000 10.2000 99.9000 ;
	    RECT 12.0000 98.2000 12.4000 99.9000 ;
	    RECT 12.0000 97.9000 13.0000 98.2000 ;
	    RECT 7.8000 97.5000 8.2000 97.9000 ;
	    RECT 9.9000 97.6000 10.2000 97.9000 ;
	    RECT 9.5000 97.3000 11.3000 97.6000 ;
	    RECT 12.6000 97.5000 13.0000 97.9000 ;
	    RECT 9.5000 97.2000 9.9000 97.3000 ;
	    RECT 10.9000 97.2000 11.3000 97.3000 ;
	    RECT 7.0000 97.0000 7.7000 97.2000 ;
	    RECT 7.0000 96.8000 8.1000 97.0000 ;
	    RECT 7.4000 96.6000 8.1000 96.8000 ;
	    RECT 7.8000 96.1000 8.1000 96.6000 ;
	    RECT 8.9000 96.5000 10.0000 96.8000 ;
	    RECT 8.9000 96.4000 9.3000 96.5000 ;
	    RECT 7.8000 95.8000 9.0000 96.1000 ;
	    RECT 5.4000 95.3000 7.5000 95.6000 ;
	    RECT 1.5000 93.7000 1.8000 95.2000 ;
	    RECT 2.2000 94.4000 2.6000 95.2000 ;
	    RECT 3.9000 93.7000 4.2000 95.2000 ;
	    RECT 4.6000 95.1000 5.0000 95.2000 ;
	    RECT 5.4000 95.1000 5.8000 95.3000 ;
	    RECT 7.1000 95.2000 7.5000 95.3000 ;
	    RECT 4.6000 94.8000 5.8000 95.1000 ;
	    RECT 4.6000 94.4000 5.0000 94.8000 ;
	    RECT 1.5000 93.4000 2.6000 93.7000 ;
	    RECT 3.9000 93.4000 5.0000 93.7000 ;
	    RECT 2.2000 91.1000 2.6000 93.4000 ;
	    RECT 4.6000 91.1000 5.0000 93.4000 ;
	    RECT 5.4000 93.6000 5.8000 94.8000 ;
	    RECT 6.3000 94.9000 6.7000 95.0000 ;
	    RECT 6.3000 94.6000 8.2000 94.9000 ;
	    RECT 7.8000 94.5000 8.2000 94.6000 ;
	    RECT 8.7000 94.2000 9.0000 95.8000 ;
	    RECT 9.7000 95.9000 10.0000 96.5000 ;
	    RECT 10.3000 96.5000 10.7000 96.6000 ;
	    RECT 12.6000 96.5000 13.0000 96.6000 ;
	    RECT 10.3000 96.2000 13.0000 96.5000 ;
	    RECT 9.7000 95.7000 12.1000 95.9000 ;
	    RECT 14.2000 95.7000 14.6000 99.9000 ;
	    RECT 9.7000 95.6000 14.6000 95.7000 ;
	    RECT 11.7000 95.5000 14.6000 95.6000 ;
	    RECT 11.8000 95.4000 14.6000 95.5000 ;
	    RECT 15.0000 95.6000 15.4000 99.9000 ;
	    RECT 17.1000 97.9000 17.7000 99.9000 ;
	    RECT 19.4000 97.9000 19.8000 99.9000 ;
	    RECT 21.6000 98.2000 22.0000 99.9000 ;
	    RECT 21.6000 97.9000 22.6000 98.2000 ;
	    RECT 17.4000 97.5000 17.8000 97.9000 ;
	    RECT 19.5000 97.6000 19.8000 97.9000 ;
	    RECT 19.1000 97.3000 20.9000 97.6000 ;
	    RECT 22.2000 97.5000 22.6000 97.9000 ;
	    RECT 19.1000 97.2000 19.5000 97.3000 ;
	    RECT 20.5000 97.2000 20.9000 97.3000 ;
	    RECT 17.0000 96.6000 17.7000 97.0000 ;
	    RECT 17.4000 96.1000 17.7000 96.6000 ;
	    RECT 18.5000 96.5000 19.6000 96.8000 ;
	    RECT 18.5000 96.4000 18.9000 96.5000 ;
	    RECT 17.4000 95.8000 18.6000 96.1000 ;
	    RECT 15.0000 95.3000 17.1000 95.6000 ;
	    RECT 11.0000 95.1000 11.4000 95.2000 ;
	    RECT 11.0000 94.8000 13.5000 95.1000 ;
	    RECT 11.8000 94.7000 12.2000 94.8000 ;
	    RECT 13.1000 94.7000 13.5000 94.8000 ;
	    RECT 12.3000 94.2000 12.7000 94.3000 ;
	    RECT 6.2000 93.6000 6.6000 94.2000 ;
	    RECT 8.7000 93.9000 14.2000 94.2000 ;
	    RECT 8.9000 93.8000 9.8000 93.9000 ;
	    RECT 5.4000 93.3000 7.3000 93.6000 ;
	    RECT 5.4000 91.1000 5.8000 93.3000 ;
	    RECT 6.9000 93.2000 7.3000 93.3000 ;
	    RECT 11.8000 92.8000 12.1000 93.9000 ;
	    RECT 13.4000 93.8000 14.2000 93.9000 ;
	    RECT 15.0000 93.6000 15.4000 95.3000 ;
	    RECT 16.7000 95.2000 17.1000 95.3000 ;
	    RECT 15.9000 94.9000 16.3000 95.0000 ;
	    RECT 15.9000 94.6000 17.8000 94.9000 ;
	    RECT 17.4000 94.5000 17.8000 94.6000 ;
	    RECT 18.3000 94.2000 18.6000 95.8000 ;
	    RECT 19.3000 95.9000 19.6000 96.5000 ;
	    RECT 19.9000 96.5000 20.3000 96.6000 ;
	    RECT 22.2000 96.5000 22.6000 96.6000 ;
	    RECT 19.9000 96.2000 22.6000 96.5000 ;
	    RECT 19.3000 95.7000 21.7000 95.9000 ;
	    RECT 23.8000 95.7000 24.2000 99.9000 ;
	    RECT 24.6000 96.2000 25.0000 99.9000 ;
	    RECT 25.4000 96.2000 25.8000 96.3000 ;
	    RECT 26.8000 96.2000 27.6000 99.9000 ;
	    RECT 24.6000 95.9000 25.8000 96.2000 ;
	    RECT 26.6000 95.9000 27.6000 96.2000 ;
	    RECT 28.7000 96.2000 29.1000 96.3000 ;
	    RECT 29.4000 96.2000 29.8000 99.9000 ;
	    RECT 28.7000 95.9000 29.8000 96.2000 ;
	    RECT 31.5000 96.2000 31.9000 99.9000 ;
	    RECT 32.2000 96.8000 32.6000 97.2000 ;
	    RECT 32.3000 96.2000 32.6000 96.8000 ;
	    RECT 34.7000 96.3000 35.1000 99.9000 ;
	    RECT 31.5000 95.9000 32.0000 96.2000 ;
	    RECT 32.3000 95.9000 33.0000 96.2000 ;
	    RECT 34.2000 95.9000 35.1000 96.3000 ;
	    RECT 35.8000 96.2000 36.2000 99.9000 ;
	    RECT 36.6000 96.2000 37.0000 96.3000 ;
	    RECT 35.8000 95.9000 37.0000 96.2000 ;
	    RECT 38.0000 95.9000 38.8000 99.9000 ;
	    RECT 39.7000 96.2000 40.1000 96.3000 ;
	    RECT 40.6000 96.2000 41.0000 99.9000 ;
	    RECT 39.7000 95.9000 41.0000 96.2000 ;
	    RECT 41.7000 96.3000 42.1000 99.9000 ;
	    RECT 45.1000 99.2000 45.5000 99.9000 ;
	    RECT 44.6000 98.8000 45.5000 99.2000 ;
	    RECT 41.7000 95.9000 42.6000 96.3000 ;
	    RECT 45.1000 96.2000 45.5000 98.8000 ;
	    RECT 45.8000 96.8000 46.2000 97.2000 ;
	    RECT 45.9000 96.2000 46.2000 96.8000 ;
	    RECT 45.1000 95.9000 45.6000 96.2000 ;
	    RECT 45.9000 96.1000 46.6000 96.2000 ;
	    RECT 48.6000 96.1000 49.0000 99.9000 ;
	    RECT 45.9000 95.9000 49.0000 96.1000 ;
	    RECT 49.4000 96.2000 49.8000 99.9000 ;
	    RECT 51.0000 96.2000 51.4000 99.9000 ;
	    RECT 49.4000 95.9000 51.4000 96.2000 ;
	    RECT 51.8000 95.9000 52.2000 99.9000 ;
	    RECT 52.6000 96.2000 53.0000 99.9000 ;
	    RECT 54.2000 96.2000 54.6000 99.9000 ;
	    RECT 52.6000 95.9000 54.6000 96.2000 ;
	    RECT 19.3000 95.6000 24.2000 95.7000 ;
	    RECT 21.3000 95.5000 24.2000 95.6000 ;
	    RECT 21.4000 95.4000 24.2000 95.5000 ;
	    RECT 26.6000 95.2000 26.9000 95.9000 ;
	    RECT 28.7000 95.6000 29.0000 95.9000 ;
	    RECT 27.3000 95.3000 29.0000 95.6000 ;
	    RECT 27.3000 95.2000 27.7000 95.3000 ;
	    RECT 20.6000 95.1000 21.0000 95.2000 ;
	    RECT 20.6000 94.8000 23.1000 95.1000 ;
	    RECT 26.2000 94.9000 26.9000 95.2000 ;
	    RECT 28.4000 94.9000 28.8000 95.0000 ;
	    RECT 26.2000 94.8000 27.1000 94.9000 ;
	    RECT 21.4000 94.7000 21.8000 94.8000 ;
	    RECT 22.7000 94.7000 23.1000 94.8000 ;
	    RECT 26.6000 94.6000 27.1000 94.8000 ;
	    RECT 21.9000 94.2000 22.3000 94.3000 ;
	    RECT 18.2000 93.9000 23.8000 94.2000 ;
	    RECT 18.2000 93.8000 18.9000 93.9000 ;
	    RECT 10.9000 92.7000 11.3000 92.8000 ;
	    RECT 7.8000 92.1000 8.2000 92.5000 ;
	    RECT 9.9000 92.4000 11.3000 92.7000 ;
	    RECT 11.8000 92.4000 12.2000 92.8000 ;
	    RECT 9.9000 92.1000 10.2000 92.4000 ;
	    RECT 12.6000 92.1000 13.0000 92.5000 ;
	    RECT 7.5000 91.8000 8.2000 92.1000 ;
	    RECT 7.5000 91.1000 8.1000 91.8000 ;
	    RECT 9.8000 91.1000 10.2000 92.1000 ;
	    RECT 12.0000 91.8000 13.0000 92.1000 ;
	    RECT 12.0000 91.1000 12.4000 91.8000 ;
	    RECT 14.2000 91.1000 14.6000 93.5000 ;
	    RECT 15.0000 93.3000 16.9000 93.6000 ;
	    RECT 15.0000 91.1000 15.4000 93.3000 ;
	    RECT 16.5000 93.2000 16.9000 93.3000 ;
	    RECT 18.2000 93.2000 18.5000 93.8000 ;
	    RECT 18.2000 92.8000 18.6000 93.2000 ;
	    RECT 21.4000 92.8000 21.7000 93.9000 ;
	    RECT 23.0000 93.8000 23.8000 93.9000 ;
	    RECT 24.6000 93.8000 25.4000 94.2000 ;
	    RECT 26.0000 93.8000 26.4000 94.2000 ;
	    RECT 26.1000 93.6000 26.4000 93.8000 ;
	    RECT 20.5000 92.7000 20.9000 92.8000 ;
	    RECT 17.4000 92.1000 17.8000 92.5000 ;
	    RECT 19.5000 92.4000 20.9000 92.7000 ;
	    RECT 21.4000 92.4000 21.8000 92.8000 ;
	    RECT 19.5000 92.1000 19.8000 92.4000 ;
	    RECT 22.2000 92.1000 22.6000 92.5000 ;
	    RECT 17.1000 91.8000 17.8000 92.1000 ;
	    RECT 17.1000 91.1000 17.7000 91.8000 ;
	    RECT 19.4000 91.1000 19.8000 92.1000 ;
	    RECT 21.6000 91.8000 22.6000 92.1000 ;
	    RECT 21.6000 91.1000 22.0000 91.8000 ;
	    RECT 23.8000 91.1000 24.2000 93.5000 ;
	    RECT 25.4000 93.4000 25.8000 93.5000 ;
	    RECT 24.6000 93.1000 25.8000 93.4000 ;
	    RECT 26.1000 93.2000 26.5000 93.6000 ;
	    RECT 24.6000 91.1000 25.0000 93.1000 ;
	    RECT 26.8000 92.9000 27.1000 94.6000 ;
	    RECT 27.5000 94.6000 28.8000 94.9000 ;
	    RECT 27.5000 94.3000 27.8000 94.6000 ;
	    RECT 31.0000 94.4000 31.4000 95.2000 ;
	    RECT 27.4000 93.9000 27.8000 94.3000 ;
	    RECT 31.7000 94.2000 32.0000 95.9000 ;
	    RECT 32.6000 95.8000 33.0000 95.9000 ;
	    RECT 33.4000 95.1000 33.8000 95.2000 ;
	    RECT 34.3000 95.1000 34.6000 95.9000 ;
	    RECT 33.4000 94.8000 34.6000 95.1000 ;
	    RECT 35.0000 94.8000 35.4000 95.6000 ;
	    RECT 38.2000 95.2000 38.5000 95.9000 ;
	    RECT 39.1000 95.2000 39.5000 95.3000 ;
	    RECT 38.2000 94.8000 38.6000 95.2000 ;
	    RECT 39.1000 94.9000 39.9000 95.2000 ;
	    RECT 39.5000 94.8000 39.9000 94.9000 ;
	    RECT 40.6000 95.1000 41.0000 95.2000 ;
	    RECT 41.4000 95.1000 41.8000 95.6000 ;
	    RECT 40.6000 94.8000 41.8000 95.1000 ;
	    RECT 34.3000 94.2000 34.6000 94.8000 ;
	    RECT 38.2000 94.2000 38.5000 94.8000 ;
	    RECT 29.0000 94.1000 29.8000 94.2000 ;
	    RECT 28.1000 93.8000 29.8000 94.1000 ;
	    RECT 30.2000 94.1000 30.6000 94.2000 ;
	    RECT 30.2000 93.8000 31.0000 94.1000 ;
	    RECT 31.7000 93.8000 33.0000 94.2000 ;
	    RECT 34.2000 93.8000 34.6000 94.2000 ;
	    RECT 35.8000 93.8000 36.6000 94.2000 ;
	    RECT 37.2000 93.8000 37.6000 94.2000 ;
	    RECT 28.1000 93.6000 28.4000 93.8000 ;
	    RECT 30.6000 93.6000 31.0000 93.8000 ;
	    RECT 27.4000 93.3000 28.4000 93.6000 ;
	    RECT 28.7000 93.4000 29.1000 93.5000 ;
	    RECT 27.4000 93.2000 28.2000 93.3000 ;
	    RECT 28.7000 93.1000 29.8000 93.4000 ;
	    RECT 30.3000 93.1000 32.1000 93.3000 ;
	    RECT 32.6000 93.1000 32.9000 93.8000 ;
	    RECT 26.8000 91.1000 27.6000 92.9000 ;
	    RECT 29.4000 91.1000 29.8000 93.1000 ;
	    RECT 30.2000 93.0000 32.2000 93.1000 ;
	    RECT 30.2000 91.1000 30.6000 93.0000 ;
	    RECT 31.8000 91.1000 32.2000 93.0000 ;
	    RECT 32.6000 91.1000 33.0000 93.1000 ;
	    RECT 33.4000 92.4000 33.8000 93.2000 ;
	    RECT 34.3000 92.1000 34.6000 93.8000 ;
	    RECT 37.3000 93.6000 37.6000 93.8000 ;
	    RECT 38.0000 93.9000 38.5000 94.2000 ;
	    RECT 38.8000 94.3000 39.2000 94.4000 ;
	    RECT 38.8000 94.2000 40.2000 94.3000 ;
	    RECT 42.2000 94.2000 42.5000 95.9000 ;
	    RECT 44.6000 94.4000 45.0000 95.2000 ;
	    RECT 45.3000 94.2000 45.6000 95.9000 ;
	    RECT 46.2000 95.8000 49.0000 95.9000 ;
	    RECT 48.7000 95.2000 49.0000 95.8000 ;
	    RECT 50.6000 95.2000 51.0000 95.4000 ;
	    RECT 51.9000 95.2000 52.2000 95.9000 ;
	    RECT 53.8000 95.2000 54.2000 95.4000 ;
	    RECT 48.6000 94.9000 49.8000 95.2000 ;
	    RECT 50.6000 94.9000 51.4000 95.2000 ;
	    RECT 48.6000 94.8000 49.0000 94.9000 ;
	    RECT 38.8000 94.0000 41.0000 94.2000 ;
	    RECT 39.9000 93.9000 41.0000 94.0000 ;
	    RECT 36.6000 93.4000 37.0000 93.5000 ;
	    RECT 34.2000 91.1000 34.6000 92.1000 ;
	    RECT 35.8000 93.1000 37.0000 93.4000 ;
	    RECT 37.3000 93.2000 37.7000 93.6000 ;
	    RECT 35.8000 91.1000 36.2000 93.1000 ;
	    RECT 38.0000 92.9000 38.3000 93.9000 ;
	    RECT 40.2000 93.8000 41.0000 93.9000 ;
	    RECT 42.2000 94.1000 42.6000 94.2000 ;
	    RECT 43.8000 94.1000 44.2000 94.2000 ;
	    RECT 42.2000 93.8000 44.6000 94.1000 ;
	    RECT 45.3000 93.8000 46.6000 94.2000 ;
	    RECT 38.6000 93.2000 39.4000 93.6000 ;
	    RECT 39.7000 93.4000 40.1000 93.5000 ;
	    RECT 39.7000 93.1000 41.0000 93.4000 ;
	    RECT 38.0000 92.2000 38.8000 92.9000 ;
	    RECT 37.4000 91.8000 38.8000 92.2000 ;
	    RECT 38.0000 91.1000 38.8000 91.8000 ;
	    RECT 40.6000 91.1000 41.0000 93.1000 ;
	    RECT 42.2000 92.1000 42.5000 93.8000 ;
	    RECT 44.2000 93.6000 44.6000 93.8000 ;
	    RECT 43.0000 92.4000 43.4000 93.2000 ;
	    RECT 43.9000 93.1000 45.7000 93.3000 ;
	    RECT 46.2000 93.1000 46.5000 93.8000 ;
	    RECT 43.8000 93.0000 45.8000 93.1000 ;
	    RECT 42.2000 91.1000 42.6000 92.1000 ;
	    RECT 43.8000 91.1000 44.2000 93.0000 ;
	    RECT 45.4000 91.1000 45.8000 93.0000 ;
	    RECT 46.2000 91.1000 46.6000 93.1000 ;
	    RECT 48.6000 92.8000 49.0000 93.2000 ;
	    RECT 49.5000 93.1000 49.8000 94.9000 ;
	    RECT 51.0000 94.8000 51.4000 94.9000 ;
	    RECT 51.8000 94.9000 53.0000 95.2000 ;
	    RECT 53.8000 94.9000 54.6000 95.2000 ;
	    RECT 51.8000 94.8000 52.2000 94.9000 ;
	    RECT 50.2000 93.8000 50.6000 94.6000 ;
	    RECT 52.7000 93.2000 53.0000 94.9000 ;
	    RECT 54.2000 94.8000 54.6000 94.9000 ;
	    RECT 53.4000 93.8000 53.8000 94.6000 ;
	    RECT 48.7000 92.4000 49.1000 92.8000 ;
	    RECT 49.4000 91.1000 49.8000 93.1000 ;
	    RECT 51.8000 92.8000 52.2000 93.2000 ;
	    RECT 51.9000 92.4000 52.3000 92.8000 ;
	    RECT 52.6000 91.1000 53.0000 93.2000 ;
	    RECT 55.0000 91.1000 55.4000 99.9000 ;
	    RECT 57.4000 97.9000 57.8000 99.9000 ;
	    RECT 57.5000 97.8000 57.8000 97.9000 ;
	    RECT 59.0000 97.9000 59.4000 99.9000 ;
	    RECT 59.0000 97.8000 59.3000 97.9000 ;
	    RECT 57.5000 97.5000 59.3000 97.8000 ;
	    RECT 58.2000 96.4000 58.6000 97.2000 ;
	    RECT 59.0000 96.2000 59.3000 97.5000 ;
	    RECT 59.8000 96.2000 60.2000 99.9000 ;
	    RECT 62.2000 96.2000 62.6000 99.9000 ;
	    RECT 63.8000 96.2000 64.2000 99.9000 ;
	    RECT 56.6000 95.4000 57.0000 96.2000 ;
	    RECT 59.0000 95.8000 59.4000 96.2000 ;
	    RECT 59.8000 95.9000 60.9000 96.2000 ;
	    RECT 62.2000 95.9000 64.2000 96.2000 ;
	    RECT 64.6000 95.9000 65.0000 99.9000 ;
	    RECT 65.8000 96.8000 66.2000 97.2000 ;
	    RECT 65.8000 96.2000 66.1000 96.8000 ;
	    RECT 66.5000 96.2000 66.9000 99.9000 ;
	    RECT 65.4000 95.9000 66.1000 96.2000 ;
	    RECT 66.4000 95.9000 66.9000 96.2000 ;
	    RECT 57.4000 94.8000 58.2000 95.2000 ;
	    RECT 59.0000 94.2000 59.3000 95.8000 ;
	    RECT 60.6000 95.6000 60.9000 95.9000 ;
	    RECT 60.6000 95.2000 61.2000 95.6000 ;
	    RECT 62.6000 95.2000 63.0000 95.4000 ;
	    RECT 64.6000 95.2000 64.9000 95.9000 ;
	    RECT 65.4000 95.8000 65.8000 95.9000 ;
	    RECT 59.8000 94.4000 60.2000 95.2000 ;
	    RECT 57.4000 93.8000 57.8000 94.2000 ;
	    RECT 58.5000 94.1000 59.3000 94.2000 ;
	    RECT 58.4000 93.9000 59.3000 94.1000 ;
	    RECT 55.8000 92.4000 56.2000 93.2000 ;
	    RECT 57.4000 93.1000 57.7000 93.8000 ;
	    RECT 58.4000 93.1000 58.8000 93.9000 ;
	    RECT 60.6000 93.7000 60.9000 95.2000 ;
	    RECT 62.2000 94.9000 63.0000 95.2000 ;
	    RECT 63.8000 94.9000 65.0000 95.2000 ;
	    RECT 62.2000 94.8000 62.6000 94.9000 ;
	    RECT 63.0000 93.8000 63.4000 94.6000 ;
	    RECT 57.4000 92.8000 58.8000 93.1000 ;
	    RECT 58.4000 91.1000 58.8000 92.8000 ;
	    RECT 59.8000 93.4000 60.9000 93.7000 ;
	    RECT 59.8000 91.1000 60.2000 93.4000 ;
	    RECT 63.8000 93.1000 64.1000 94.9000 ;
	    RECT 64.6000 94.8000 65.0000 94.9000 ;
	    RECT 66.4000 94.2000 66.7000 95.9000 ;
	    RECT 67.0000 95.1000 67.4000 95.2000 ;
	    RECT 67.8000 95.1000 68.2000 95.2000 ;
	    RECT 67.0000 94.8000 68.2000 95.1000 ;
	    RECT 67.0000 94.4000 67.4000 94.8000 ;
	    RECT 65.4000 93.8000 66.7000 94.2000 ;
	    RECT 67.8000 94.1000 68.2000 94.2000 ;
	    RECT 67.4000 93.8000 68.2000 94.1000 ;
	    RECT 64.6000 93.1000 65.0000 93.2000 ;
	    RECT 65.5000 93.1000 65.8000 93.8000 ;
	    RECT 67.4000 93.6000 67.8000 93.8000 ;
	    RECT 66.3000 93.1000 68.1000 93.3000 ;
	    RECT 63.8000 91.1000 64.2000 93.1000 ;
	    RECT 64.6000 92.8000 65.8000 93.1000 ;
	    RECT 64.5000 92.4000 64.9000 92.8000 ;
	    RECT 65.4000 91.1000 65.8000 92.8000 ;
	    RECT 66.2000 93.0000 68.2000 93.1000 ;
	    RECT 66.2000 91.1000 66.6000 93.0000 ;
	    RECT 67.8000 91.1000 68.2000 93.0000 ;
	    RECT 68.6000 92.4000 69.0000 93.2000 ;
	    RECT 69.4000 93.1000 69.8000 99.9000 ;
	    RECT 71.5000 96.3000 71.9000 99.9000 ;
	    RECT 71.0000 95.9000 71.9000 96.3000 ;
	    RECT 70.2000 95.1000 70.6000 95.2000 ;
	    RECT 71.1000 95.1000 71.4000 95.9000 ;
	    RECT 72.6000 95.7000 73.0000 99.9000 ;
	    RECT 74.8000 98.2000 75.2000 99.9000 ;
	    RECT 74.2000 97.9000 75.2000 98.2000 ;
	    RECT 77.0000 97.9000 77.4000 99.9000 ;
	    RECT 79.1000 97.9000 79.7000 99.9000 ;
	    RECT 74.2000 97.5000 74.6000 97.9000 ;
	    RECT 77.0000 97.6000 77.3000 97.9000 ;
	    RECT 75.9000 97.3000 77.7000 97.6000 ;
	    RECT 79.0000 97.5000 79.4000 97.9000 ;
	    RECT 75.9000 97.2000 76.3000 97.3000 ;
	    RECT 77.3000 97.2000 77.7000 97.3000 ;
	    RECT 74.2000 96.5000 74.6000 96.6000 ;
	    RECT 76.5000 96.5000 76.9000 96.6000 ;
	    RECT 74.2000 96.2000 76.9000 96.5000 ;
	    RECT 77.2000 96.5000 78.3000 96.8000 ;
	    RECT 77.2000 95.9000 77.5000 96.5000 ;
	    RECT 77.9000 96.4000 78.3000 96.5000 ;
	    RECT 79.1000 96.6000 79.8000 97.0000 ;
	    RECT 79.1000 96.1000 79.4000 96.6000 ;
	    RECT 75.1000 95.7000 77.5000 95.9000 ;
	    RECT 72.6000 95.6000 77.5000 95.7000 ;
	    RECT 78.2000 95.8000 79.4000 96.1000 ;
	    RECT 70.2000 94.8000 71.4000 95.1000 ;
	    RECT 71.8000 94.8000 72.2000 95.6000 ;
	    RECT 72.6000 95.5000 75.5000 95.6000 ;
	    RECT 72.6000 95.4000 75.4000 95.5000 ;
	    RECT 78.2000 95.2000 78.5000 95.8000 ;
	    RECT 81.4000 95.6000 81.8000 99.9000 ;
	    RECT 82.2000 96.2000 82.6000 99.9000 ;
	    RECT 82.2000 95.9000 83.3000 96.2000 ;
	    RECT 83.8000 95.9000 84.2000 99.9000 ;
	    RECT 79.7000 95.3000 81.8000 95.6000 ;
	    RECT 79.7000 95.2000 80.1000 95.3000 ;
	    RECT 75.8000 95.1000 76.2000 95.2000 ;
	    RECT 73.7000 94.8000 76.2000 95.1000 ;
	    RECT 78.2000 94.8000 78.6000 95.2000 ;
	    RECT 80.5000 94.9000 80.9000 95.0000 ;
	    RECT 71.1000 94.2000 71.4000 94.8000 ;
	    RECT 73.7000 94.7000 74.1000 94.8000 ;
	    RECT 75.0000 94.7000 75.4000 94.8000 ;
	    RECT 74.5000 94.2000 74.9000 94.3000 ;
	    RECT 78.2000 94.2000 78.5000 94.8000 ;
	    RECT 79.0000 94.6000 80.9000 94.9000 ;
	    RECT 79.0000 94.5000 79.4000 94.6000 ;
	    RECT 71.0000 93.8000 71.4000 94.2000 ;
	    RECT 73.0000 93.9000 78.5000 94.2000 ;
	    RECT 73.0000 93.8000 73.8000 93.9000 ;
	    RECT 70.2000 93.1000 70.6000 93.2000 ;
	    RECT 69.4000 92.8000 70.6000 93.1000 ;
	    RECT 69.4000 91.1000 69.8000 92.8000 ;
	    RECT 70.2000 92.4000 70.6000 92.8000 ;
	    RECT 71.1000 92.1000 71.4000 93.8000 ;
	    RECT 71.0000 91.1000 71.4000 92.1000 ;
	    RECT 72.6000 91.1000 73.0000 93.5000 ;
	    RECT 75.1000 92.8000 75.4000 93.9000 ;
	    RECT 77.9000 93.8000 78.3000 93.9000 ;
	    RECT 81.4000 93.6000 81.8000 95.3000 ;
	    RECT 83.0000 95.6000 83.3000 95.9000 ;
	    RECT 83.0000 95.2000 83.6000 95.6000 ;
	    RECT 82.2000 94.4000 82.6000 95.2000 ;
	    RECT 83.0000 93.7000 83.3000 95.2000 ;
	    RECT 83.9000 94.8000 84.2000 95.9000 ;
	    RECT 79.9000 93.3000 81.8000 93.6000 ;
	    RECT 79.9000 93.2000 80.3000 93.3000 ;
	    RECT 74.2000 92.1000 74.6000 92.5000 ;
	    RECT 75.0000 92.4000 75.4000 92.8000 ;
	    RECT 75.9000 92.7000 76.3000 92.8000 ;
	    RECT 75.9000 92.4000 77.3000 92.7000 ;
	    RECT 77.0000 92.1000 77.3000 92.4000 ;
	    RECT 79.0000 92.1000 79.4000 92.5000 ;
	    RECT 74.2000 91.8000 75.2000 92.1000 ;
	    RECT 74.8000 91.1000 75.2000 91.8000 ;
	    RECT 77.0000 91.1000 77.4000 92.1000 ;
	    RECT 79.0000 91.8000 79.7000 92.1000 ;
	    RECT 79.1000 91.1000 79.7000 91.8000 ;
	    RECT 81.4000 91.1000 81.8000 93.3000 ;
	    RECT 82.2000 93.4000 83.3000 93.7000 ;
	    RECT 82.2000 91.1000 82.6000 93.4000 ;
	    RECT 83.8000 91.1000 84.2000 94.8000 ;
	    RECT 84.6000 95.9000 85.0000 99.9000 ;
	    RECT 86.2000 96.2000 86.6000 99.9000 ;
	    RECT 88.9000 99.2000 89.3000 99.9000 ;
	    RECT 88.9000 98.8000 89.8000 99.2000 ;
	    RECT 88.9000 96.4000 89.3000 98.8000 ;
	    RECT 91.0000 97.5000 91.4000 99.5000 ;
	    RECT 85.5000 95.9000 86.6000 96.2000 ;
	    RECT 88.5000 96.1000 89.3000 96.4000 ;
	    RECT 84.6000 94.8000 84.9000 95.9000 ;
	    RECT 85.5000 95.6000 85.8000 95.9000 ;
	    RECT 85.2000 95.2000 85.8000 95.6000 ;
	    RECT 84.6000 91.1000 85.0000 94.8000 ;
	    RECT 85.5000 93.7000 85.8000 95.2000 ;
	    RECT 86.2000 94.4000 86.6000 95.2000 ;
	    RECT 87.8000 94.8000 88.2000 95.6000 ;
	    RECT 88.5000 94.2000 88.8000 96.1000 ;
	    RECT 91.1000 95.8000 91.4000 97.5000 ;
	    RECT 91.8000 96.2000 92.2000 99.9000 ;
	    RECT 91.8000 95.9000 92.9000 96.2000 ;
	    RECT 93.4000 95.9000 93.8000 99.9000 ;
	    RECT 95.5000 99.2000 95.9000 99.9000 ;
	    RECT 95.0000 98.8000 95.9000 99.2000 ;
	    RECT 95.5000 96.3000 95.9000 98.8000 ;
	    RECT 95.0000 95.9000 95.9000 96.3000 ;
	    RECT 89.5000 95.5000 91.4000 95.8000 ;
	    RECT 92.6000 95.6000 92.9000 95.9000 ;
	    RECT 89.5000 94.5000 89.8000 95.5000 ;
	    RECT 92.6000 95.2000 93.2000 95.6000 ;
	    RECT 87.8000 93.8000 88.8000 94.2000 ;
	    RECT 89.1000 94.1000 89.8000 94.5000 ;
	    RECT 90.2000 94.4000 90.6000 95.2000 ;
	    RECT 91.0000 94.4000 91.4000 95.2000 ;
	    RECT 91.8000 94.4000 92.2000 95.2000 ;
	    RECT 85.5000 93.4000 86.6000 93.7000 ;
	    RECT 86.2000 91.1000 86.6000 93.4000 ;
	    RECT 88.5000 93.5000 88.8000 93.8000 ;
	    RECT 89.3000 93.9000 89.8000 94.1000 ;
	    RECT 89.3000 93.6000 91.4000 93.9000 ;
	    RECT 92.6000 93.7000 92.9000 95.2000 ;
	    RECT 93.5000 94.8000 93.8000 95.9000 ;
	    RECT 88.5000 93.3000 88.9000 93.5000 ;
	    RECT 88.5000 93.0000 89.3000 93.3000 ;
	    RECT 88.9000 91.5000 89.3000 93.0000 ;
	    RECT 91.1000 92.5000 91.4000 93.6000 ;
	    RECT 91.0000 91.5000 91.4000 92.5000 ;
	    RECT 91.8000 93.4000 92.9000 93.7000 ;
	    RECT 91.8000 91.1000 92.2000 93.4000 ;
	    RECT 93.4000 91.1000 93.8000 94.8000 ;
	    RECT 95.1000 94.2000 95.4000 95.9000 ;
	    RECT 95.8000 95.1000 96.2000 95.6000 ;
	    RECT 96.6000 95.1000 97.0000 99.9000 ;
	    RECT 101.4000 96.2000 101.8000 99.9000 ;
	    RECT 100.7000 95.9000 101.8000 96.2000 ;
	    RECT 100.7000 95.6000 101.0000 95.9000 ;
	    RECT 100.4000 95.2000 101.0000 95.6000 ;
	    RECT 102.2000 95.6000 102.6000 99.9000 ;
	    RECT 104.3000 97.9000 104.9000 99.9000 ;
	    RECT 106.6000 97.9000 107.0000 99.9000 ;
	    RECT 108.8000 98.2000 109.2000 99.9000 ;
	    RECT 108.8000 97.9000 109.8000 98.2000 ;
	    RECT 104.6000 97.5000 105.0000 97.9000 ;
	    RECT 106.7000 97.6000 107.0000 97.9000 ;
	    RECT 106.3000 97.3000 108.1000 97.6000 ;
	    RECT 109.4000 97.5000 109.8000 97.9000 ;
	    RECT 106.3000 97.2000 106.7000 97.3000 ;
	    RECT 107.7000 97.2000 108.1000 97.3000 ;
	    RECT 104.2000 96.6000 104.9000 97.0000 ;
	    RECT 104.6000 96.1000 104.9000 96.6000 ;
	    RECT 105.7000 96.5000 106.8000 96.8000 ;
	    RECT 105.7000 96.4000 106.1000 96.5000 ;
	    RECT 104.6000 95.8000 105.8000 96.1000 ;
	    RECT 102.2000 95.3000 104.3000 95.6000 ;
	    RECT 95.8000 94.8000 97.0000 95.1000 ;
	    RECT 95.0000 93.8000 95.4000 94.2000 ;
	    RECT 94.2000 92.4000 94.6000 93.2000 ;
	    RECT 95.1000 92.2000 95.4000 93.8000 ;
	    RECT 95.0000 91.1000 95.4000 92.2000 ;
	    RECT 96.6000 91.1000 97.0000 94.8000 ;
	    RECT 97.4000 93.4000 97.8000 94.2000 ;
	    RECT 100.7000 93.7000 101.0000 95.2000 ;
	    RECT 101.4000 95.1000 101.8000 95.2000 ;
	    RECT 102.2000 95.1000 102.6000 95.3000 ;
	    RECT 103.9000 95.2000 104.3000 95.3000 ;
	    RECT 105.5000 95.2000 105.8000 95.8000 ;
	    RECT 106.5000 95.9000 106.8000 96.5000 ;
	    RECT 107.1000 96.5000 107.5000 96.6000 ;
	    RECT 109.4000 96.5000 109.8000 96.6000 ;
	    RECT 107.1000 96.2000 109.8000 96.5000 ;
	    RECT 106.5000 95.7000 108.9000 95.9000 ;
	    RECT 111.0000 95.7000 111.4000 99.9000 ;
	    RECT 112.2000 96.8000 112.6000 97.2000 ;
	    RECT 112.2000 96.2000 112.5000 96.8000 ;
	    RECT 112.9000 96.2000 113.3000 99.9000 ;
	    RECT 115.4000 96.8000 115.8000 97.2000 ;
	    RECT 115.4000 96.2000 115.7000 96.8000 ;
	    RECT 116.1000 96.2000 116.5000 99.9000 ;
	    RECT 119.0000 97.9000 119.4000 99.9000 ;
	    RECT 111.8000 95.9000 112.5000 96.2000 ;
	    RECT 112.8000 95.9000 113.3000 96.2000 ;
	    RECT 115.0000 95.9000 115.7000 96.2000 ;
	    RECT 111.8000 95.8000 112.2000 95.9000 ;
	    RECT 106.5000 95.6000 111.4000 95.7000 ;
	    RECT 108.5000 95.5000 111.4000 95.6000 ;
	    RECT 108.6000 95.4000 111.4000 95.5000 ;
	    RECT 101.4000 94.8000 102.6000 95.1000 ;
	    RECT 101.4000 94.4000 101.8000 94.8000 ;
	    RECT 100.7000 93.4000 101.8000 93.7000 ;
	    RECT 101.4000 91.1000 101.8000 93.4000 ;
	    RECT 102.2000 93.6000 102.6000 94.8000 ;
	    RECT 103.1000 94.9000 103.5000 95.0000 ;
	    RECT 103.1000 94.6000 105.0000 94.9000 ;
	    RECT 105.4000 94.8000 105.8000 95.2000 ;
	    RECT 107.8000 95.1000 108.2000 95.2000 ;
	    RECT 107.8000 94.8000 110.3000 95.1000 ;
	    RECT 104.6000 94.5000 105.0000 94.6000 ;
	    RECT 105.5000 94.2000 105.8000 94.8000 ;
	    RECT 108.6000 94.7000 109.0000 94.8000 ;
	    RECT 109.9000 94.7000 110.3000 94.8000 ;
	    RECT 109.1000 94.2000 109.5000 94.3000 ;
	    RECT 112.8000 94.2000 113.1000 95.9000 ;
	    RECT 115.0000 95.8000 115.4000 95.9000 ;
	    RECT 116.0000 95.8000 117.0000 96.2000 ;
	    RECT 119.1000 95.8000 119.4000 97.9000 ;
	    RECT 120.6000 95.9000 121.0000 99.9000 ;
	    RECT 122.7000 96.2000 123.1000 99.9000 ;
	    RECT 125.9000 97.2000 126.3000 99.9000 ;
	    RECT 123.4000 96.8000 123.8000 97.2000 ;
	    RECT 125.4000 96.8000 126.3000 97.2000 ;
	    RECT 126.6000 96.8000 127.0000 97.2000 ;
	    RECT 123.5000 96.2000 123.8000 96.8000 ;
	    RECT 125.9000 96.2000 126.3000 96.8000 ;
	    RECT 126.7000 96.2000 127.0000 96.8000 ;
	    RECT 122.7000 95.9000 123.2000 96.2000 ;
	    RECT 123.5000 95.9000 124.2000 96.2000 ;
	    RECT 125.9000 95.9000 126.4000 96.2000 ;
	    RECT 126.7000 95.9000 127.4000 96.2000 ;
	    RECT 113.4000 94.4000 113.8000 95.2000 ;
	    RECT 116.0000 94.2000 116.3000 95.8000 ;
	    RECT 119.1000 95.5000 120.3000 95.8000 ;
	    RECT 116.6000 95.1000 117.0000 95.2000 ;
	    RECT 117.4000 95.1000 117.8000 95.2000 ;
	    RECT 116.6000 94.8000 117.8000 95.1000 ;
	    RECT 119.0000 94.8000 119.4000 95.2000 ;
	    RECT 116.6000 94.4000 117.0000 94.8000 ;
	    RECT 105.5000 93.9000 111.0000 94.2000 ;
	    RECT 105.7000 93.8000 106.1000 93.9000 ;
	    RECT 102.2000 93.3000 104.2000 93.6000 ;
	    RECT 102.2000 91.1000 102.6000 93.3000 ;
	    RECT 103.7000 93.2000 104.2000 93.3000 ;
	    RECT 103.8000 92.8000 104.2000 93.2000 ;
	    RECT 108.6000 92.8000 108.9000 93.9000 ;
	    RECT 110.2000 93.8000 111.0000 93.9000 ;
	    RECT 111.8000 93.8000 113.1000 94.2000 ;
	    RECT 114.2000 94.1000 114.6000 94.2000 ;
	    RECT 113.8000 93.8000 114.6000 94.1000 ;
	    RECT 115.0000 93.8000 116.3000 94.2000 ;
	    RECT 117.4000 94.1000 117.8000 94.2000 ;
	    RECT 118.2000 94.1000 118.6000 94.6000 ;
	    RECT 119.1000 94.4000 119.4000 94.8000 ;
	    RECT 119.1000 94.1000 119.6000 94.4000 ;
	    RECT 117.0000 93.8000 118.6000 94.1000 ;
	    RECT 119.2000 94.0000 119.6000 94.1000 ;
	    RECT 120.0000 93.8000 120.3000 95.5000 ;
	    RECT 120.7000 95.2000 121.0000 95.9000 ;
	    RECT 120.6000 95.1000 121.0000 95.2000 ;
	    RECT 120.6000 94.8000 121.7000 95.1000 ;
	    RECT 107.7000 92.7000 108.1000 92.8000 ;
	    RECT 104.6000 92.1000 105.0000 92.5000 ;
	    RECT 106.7000 92.4000 108.1000 92.7000 ;
	    RECT 108.6000 92.4000 109.0000 92.8000 ;
	    RECT 106.7000 92.1000 107.0000 92.4000 ;
	    RECT 109.4000 92.1000 109.8000 92.5000 ;
	    RECT 104.3000 91.8000 105.0000 92.1000 ;
	    RECT 104.3000 91.1000 104.9000 91.8000 ;
	    RECT 106.6000 91.1000 107.0000 92.1000 ;
	    RECT 108.8000 91.8000 109.8000 92.1000 ;
	    RECT 108.8000 91.1000 109.2000 91.8000 ;
	    RECT 111.0000 91.1000 111.4000 93.5000 ;
	    RECT 111.9000 93.1000 112.2000 93.8000 ;
	    RECT 113.8000 93.6000 114.2000 93.8000 ;
	    RECT 112.7000 93.1000 114.5000 93.3000 ;
	    RECT 115.1000 93.1000 115.4000 93.8000 ;
	    RECT 117.0000 93.6000 117.4000 93.8000 ;
	    RECT 120.0000 93.7000 120.4000 93.8000 ;
	    RECT 118.9000 93.5000 120.4000 93.7000 ;
	    RECT 118.3000 93.4000 120.4000 93.5000 ;
	    RECT 115.9000 93.1000 117.7000 93.3000 ;
	    RECT 118.3000 93.2000 119.2000 93.4000 ;
	    RECT 118.3000 93.1000 118.6000 93.2000 ;
	    RECT 120.7000 93.1000 121.0000 94.8000 ;
	    RECT 121.4000 94.2000 121.7000 94.8000 ;
	    RECT 122.2000 94.4000 122.6000 95.2000 ;
	    RECT 122.9000 94.2000 123.2000 95.9000 ;
	    RECT 123.8000 95.8000 124.2000 95.9000 ;
	    RECT 125.4000 94.4000 125.8000 95.2000 ;
	    RECT 126.1000 94.2000 126.4000 95.9000 ;
	    RECT 127.0000 95.8000 127.4000 95.9000 ;
	    RECT 127.8000 95.7000 128.2000 99.9000 ;
	    RECT 130.0000 98.2000 130.4000 99.9000 ;
	    RECT 129.4000 97.9000 130.4000 98.2000 ;
	    RECT 132.2000 97.9000 132.6000 99.9000 ;
	    RECT 134.3000 97.9000 134.9000 99.9000 ;
	    RECT 129.4000 97.5000 129.8000 97.9000 ;
	    RECT 132.2000 97.6000 132.5000 97.9000 ;
	    RECT 131.1000 97.3000 132.9000 97.6000 ;
	    RECT 134.2000 97.5000 134.6000 97.9000 ;
	    RECT 131.1000 97.2000 131.5000 97.3000 ;
	    RECT 132.5000 97.2000 132.9000 97.3000 ;
	    RECT 129.4000 96.5000 129.8000 96.6000 ;
	    RECT 131.7000 96.5000 132.1000 96.6000 ;
	    RECT 129.4000 96.2000 132.1000 96.5000 ;
	    RECT 132.4000 96.5000 133.5000 96.8000 ;
	    RECT 132.4000 95.9000 132.7000 96.5000 ;
	    RECT 133.1000 96.4000 133.5000 96.5000 ;
	    RECT 134.3000 96.6000 135.0000 97.0000 ;
	    RECT 134.3000 96.1000 134.6000 96.6000 ;
	    RECT 130.3000 95.7000 132.7000 95.9000 ;
	    RECT 127.8000 95.6000 132.7000 95.7000 ;
	    RECT 133.4000 95.8000 134.6000 96.1000 ;
	    RECT 127.8000 95.5000 130.7000 95.6000 ;
	    RECT 127.8000 95.4000 130.6000 95.5000 ;
	    RECT 133.4000 95.2000 133.7000 95.8000 ;
	    RECT 136.6000 95.6000 137.0000 99.9000 ;
	    RECT 137.4000 95.9000 137.8000 99.9000 ;
	    RECT 138.2000 96.2000 138.6000 99.9000 ;
	    RECT 139.8000 96.2000 140.2000 99.9000 ;
	    RECT 138.2000 95.9000 140.2000 96.2000 ;
	    RECT 140.6000 96.2000 141.0000 99.9000 ;
	    RECT 140.6000 95.9000 141.7000 96.2000 ;
	    RECT 134.9000 95.3000 137.0000 95.6000 ;
	    RECT 134.9000 95.2000 135.3000 95.3000 ;
	    RECT 131.0000 95.1000 131.4000 95.2000 ;
	    RECT 128.9000 94.8000 131.4000 95.1000 ;
	    RECT 133.4000 94.8000 133.8000 95.2000 ;
	    RECT 135.7000 94.9000 136.1000 95.0000 ;
	    RECT 128.9000 94.7000 129.3000 94.8000 ;
	    RECT 130.2000 94.7000 130.6000 94.8000 ;
	    RECT 129.7000 94.2000 130.1000 94.3000 ;
	    RECT 133.4000 94.2000 133.7000 94.8000 ;
	    RECT 134.2000 94.6000 136.1000 94.9000 ;
	    RECT 134.2000 94.5000 134.6000 94.6000 ;
	    RECT 121.4000 94.1000 121.8000 94.2000 ;
	    RECT 121.4000 93.8000 122.2000 94.1000 ;
	    RECT 122.9000 93.8000 124.2000 94.2000 ;
	    RECT 124.6000 94.1000 125.0000 94.2000 ;
	    RECT 124.6000 93.8000 125.4000 94.1000 ;
	    RECT 126.1000 93.8000 127.4000 94.2000 ;
	    RECT 128.2000 93.9000 133.7000 94.2000 ;
	    RECT 128.2000 93.8000 129.0000 93.9000 ;
	    RECT 121.8000 93.6000 122.2000 93.8000 ;
	    RECT 121.5000 93.1000 123.3000 93.3000 ;
	    RECT 123.8000 93.1000 124.1000 93.8000 ;
	    RECT 125.0000 93.6000 125.4000 93.8000 ;
	    RECT 124.7000 93.1000 126.5000 93.3000 ;
	    RECT 127.0000 93.1000 127.3000 93.8000 ;
	    RECT 111.8000 91.1000 112.2000 93.1000 ;
	    RECT 112.6000 93.0000 114.6000 93.1000 ;
	    RECT 112.6000 91.1000 113.0000 93.0000 ;
	    RECT 114.2000 91.1000 114.6000 93.0000 ;
	    RECT 115.0000 91.1000 115.4000 93.1000 ;
	    RECT 115.8000 93.0000 117.8000 93.1000 ;
	    RECT 115.8000 91.1000 116.2000 93.0000 ;
	    RECT 117.4000 91.1000 117.8000 93.0000 ;
	    RECT 118.2000 91.1000 118.6000 93.1000 ;
	    RECT 120.3000 92.6000 121.0000 93.1000 ;
	    RECT 121.4000 93.0000 123.4000 93.1000 ;
	    RECT 120.3000 91.1000 120.7000 92.6000 ;
	    RECT 121.4000 91.1000 121.8000 93.0000 ;
	    RECT 123.0000 91.1000 123.4000 93.0000 ;
	    RECT 123.8000 91.1000 124.2000 93.1000 ;
	    RECT 124.6000 93.0000 126.6000 93.1000 ;
	    RECT 124.6000 91.1000 125.0000 93.0000 ;
	    RECT 126.2000 91.1000 126.6000 93.0000 ;
	    RECT 127.0000 91.1000 127.4000 93.1000 ;
	    RECT 127.8000 91.1000 128.2000 93.5000 ;
	    RECT 130.3000 92.8000 130.6000 93.9000 ;
	    RECT 133.1000 93.8000 133.5000 93.9000 ;
	    RECT 136.6000 93.6000 137.0000 95.3000 ;
	    RECT 137.5000 95.2000 137.8000 95.9000 ;
	    RECT 141.4000 95.6000 141.7000 95.9000 ;
	    RECT 139.4000 95.2000 139.8000 95.4000 ;
	    RECT 141.4000 95.2000 142.0000 95.6000 ;
	    RECT 137.4000 94.9000 138.6000 95.2000 ;
	    RECT 139.4000 94.9000 140.2000 95.2000 ;
	    RECT 137.4000 94.8000 137.8000 94.9000 ;
	    RECT 137.4000 94.1000 137.8000 94.2000 ;
	    RECT 138.3000 94.1000 138.6000 94.9000 ;
	    RECT 139.8000 94.8000 140.2000 94.9000 ;
	    RECT 137.4000 93.8000 138.6000 94.1000 ;
	    RECT 139.0000 93.8000 139.4000 94.6000 ;
	    RECT 140.6000 94.4000 141.0000 95.2000 ;
	    RECT 135.1000 93.3000 137.0000 93.6000 ;
	    RECT 135.1000 93.2000 135.5000 93.3000 ;
	    RECT 129.4000 92.1000 129.8000 92.5000 ;
	    RECT 130.2000 92.4000 130.6000 92.8000 ;
	    RECT 131.1000 92.7000 131.5000 92.8000 ;
	    RECT 131.1000 92.4000 132.5000 92.7000 ;
	    RECT 132.2000 92.1000 132.5000 92.4000 ;
	    RECT 134.2000 92.1000 134.6000 92.5000 ;
	    RECT 129.4000 91.8000 130.4000 92.1000 ;
	    RECT 130.0000 91.1000 130.4000 91.8000 ;
	    RECT 132.2000 91.1000 132.6000 92.1000 ;
	    RECT 134.2000 91.8000 134.9000 92.1000 ;
	    RECT 134.3000 91.1000 134.9000 91.8000 ;
	    RECT 136.6000 91.1000 137.0000 93.3000 ;
	    RECT 137.4000 92.8000 137.8000 93.2000 ;
	    RECT 138.3000 93.1000 138.6000 93.8000 ;
	    RECT 141.4000 93.7000 141.7000 95.2000 ;
	    RECT 137.5000 92.4000 137.9000 92.8000 ;
	    RECT 138.2000 91.1000 138.6000 93.1000 ;
	    RECT 140.6000 93.4000 141.7000 93.7000 ;
	    RECT 140.6000 91.1000 141.0000 93.4000 ;
	    RECT 143.0000 91.1000 143.4000 99.9000 ;
	    RECT 144.6000 96.2000 145.0000 99.9000 ;
	    RECT 144.6000 95.9000 145.7000 96.2000 ;
	    RECT 145.4000 95.6000 145.7000 95.9000 ;
	    RECT 145.4000 95.2000 146.0000 95.6000 ;
	    RECT 144.6000 94.4000 145.0000 95.2000 ;
	    RECT 145.4000 93.7000 145.7000 95.2000 ;
	    RECT 144.6000 93.4000 145.7000 93.7000 ;
	    RECT 144.6000 91.1000 145.0000 93.4000 ;
	    RECT 2.2000 87.6000 2.6000 89.9000 ;
	    RECT 1.5000 87.3000 2.6000 87.6000 ;
	    RECT 3.0000 87.7000 3.4000 89.9000 ;
	    RECT 5.1000 89.2000 5.7000 89.9000 ;
	    RECT 5.1000 88.9000 5.8000 89.2000 ;
	    RECT 7.4000 88.9000 7.8000 89.9000 ;
	    RECT 9.6000 89.2000 10.0000 89.9000 ;
	    RECT 9.6000 88.9000 10.6000 89.2000 ;
	    RECT 5.4000 88.5000 5.8000 88.9000 ;
	    RECT 7.5000 88.6000 7.8000 88.9000 ;
	    RECT 7.5000 88.3000 8.9000 88.6000 ;
	    RECT 8.5000 88.2000 8.9000 88.3000 ;
	    RECT 4.6000 87.8000 5.0000 88.2000 ;
	    RECT 4.5000 87.7000 5.0000 87.8000 ;
	    RECT 3.0000 87.4000 5.0000 87.7000 ;
	    RECT 9.4000 87.8000 9.8000 88.6000 ;
	    RECT 10.2000 88.5000 10.6000 88.9000 ;
	    RECT 1.5000 85.8000 1.8000 87.3000 ;
	    RECT 2.2000 86.1000 2.6000 86.6000 ;
	    RECT 3.0000 86.1000 3.4000 87.4000 ;
	    RECT 6.5000 87.1000 6.9000 87.2000 ;
	    RECT 9.4000 87.1000 9.7000 87.8000 ;
	    RECT 11.8000 87.5000 12.2000 89.9000 ;
	    RECT 12.6000 87.9000 13.0000 89.9000 ;
	    RECT 14.8000 89.2000 15.6000 89.9000 ;
	    RECT 14.2000 88.8000 15.6000 89.2000 ;
	    RECT 14.8000 88.1000 15.6000 88.8000 ;
	    RECT 12.6000 87.6000 13.8000 87.9000 ;
	    RECT 13.4000 87.5000 13.8000 87.6000 ;
	    RECT 14.1000 87.4000 14.5000 87.8000 ;
	    RECT 14.1000 87.2000 14.4000 87.4000 ;
	    RECT 11.0000 87.1000 11.8000 87.2000 ;
	    RECT 6.3000 86.8000 11.8000 87.1000 ;
	    RECT 12.6000 86.8000 13.4000 87.2000 ;
	    RECT 14.0000 86.8000 14.4000 87.2000 ;
	    RECT 5.4000 86.4000 5.8000 86.5000 ;
	    RECT 2.2000 85.8000 3.4000 86.1000 ;
	    RECT 3.9000 86.1000 5.8000 86.4000 ;
	    RECT 3.9000 86.0000 4.3000 86.1000 ;
	    RECT 1.2000 85.4000 1.8000 85.8000 ;
	    RECT 1.5000 85.1000 1.8000 85.4000 ;
	    RECT 3.0000 85.7000 3.4000 85.8000 ;
	    RECT 4.7000 85.7000 5.1000 85.8000 ;
	    RECT 3.0000 85.4000 5.1000 85.7000 ;
	    RECT 1.5000 84.8000 2.6000 85.1000 ;
	    RECT 2.2000 81.1000 2.6000 84.8000 ;
	    RECT 3.0000 81.1000 3.4000 85.4000 ;
	    RECT 6.3000 85.2000 6.6000 86.8000 ;
	    RECT 9.9000 86.7000 10.3000 86.8000 ;
	    RECT 14.8000 86.4000 15.1000 88.1000 ;
	    RECT 17.4000 87.9000 17.8000 89.9000 ;
	    RECT 18.2000 88.0000 18.6000 89.9000 ;
	    RECT 19.8000 88.0000 20.2000 89.9000 ;
	    RECT 18.2000 87.9000 20.2000 88.0000 ;
	    RECT 20.6000 87.9000 21.0000 89.9000 ;
	    RECT 15.4000 87.7000 16.2000 87.8000 ;
	    RECT 15.4000 87.4000 16.4000 87.7000 ;
	    RECT 16.7000 87.6000 17.8000 87.9000 ;
	    RECT 18.3000 87.7000 20.1000 87.9000 ;
	    RECT 16.7000 87.5000 17.1000 87.6000 ;
	    RECT 16.1000 87.2000 16.4000 87.4000 ;
	    RECT 18.6000 87.2000 19.0000 87.4000 ;
	    RECT 20.6000 87.2000 20.9000 87.9000 ;
	    RECT 21.4000 87.6000 21.8000 89.9000 ;
	    RECT 23.0000 88.2000 23.4000 89.9000 ;
	    RECT 23.0000 87.9000 23.5000 88.2000 ;
	    RECT 21.4000 87.3000 22.7000 87.6000 ;
	    RECT 15.4000 86.7000 15.8000 87.1000 ;
	    RECT 16.1000 86.9000 17.8000 87.2000 ;
	    RECT 17.0000 86.8000 17.8000 86.9000 ;
	    RECT 18.2000 86.9000 19.0000 87.2000 ;
	    RECT 18.2000 86.8000 18.6000 86.9000 ;
	    RECT 19.7000 86.8000 21.0000 87.2000 ;
	    RECT 9.4000 86.2000 9.8000 86.3000 ;
	    RECT 10.7000 86.2000 11.1000 86.3000 ;
	    RECT 14.6000 86.2000 15.1000 86.4000 ;
	    RECT 8.6000 85.9000 11.1000 86.2000 ;
	    RECT 14.2000 86.1000 15.1000 86.2000 ;
	    RECT 15.5000 86.4000 15.8000 86.7000 ;
	    RECT 15.5000 86.1000 16.8000 86.4000 ;
	    RECT 8.6000 85.8000 9.0000 85.9000 ;
	    RECT 14.2000 85.8000 14.9000 86.1000 ;
	    RECT 16.4000 86.0000 16.8000 86.1000 ;
	    RECT 19.0000 85.8000 19.4000 86.6000 ;
	    RECT 9.4000 85.5000 12.2000 85.6000 ;
	    RECT 9.3000 85.4000 12.2000 85.5000 ;
	    RECT 5.4000 84.9000 6.6000 85.2000 ;
	    RECT 7.3000 85.3000 12.2000 85.4000 ;
	    RECT 7.3000 85.1000 9.7000 85.3000 ;
	    RECT 5.4000 84.4000 5.7000 84.9000 ;
	    RECT 5.0000 84.0000 5.7000 84.4000 ;
	    RECT 6.5000 84.5000 6.9000 84.6000 ;
	    RECT 7.3000 84.5000 7.6000 85.1000 ;
	    RECT 6.5000 84.2000 7.6000 84.5000 ;
	    RECT 7.9000 84.5000 10.6000 84.8000 ;
	    RECT 7.9000 84.4000 8.3000 84.5000 ;
	    RECT 10.2000 84.4000 10.6000 84.5000 ;
	    RECT 7.1000 83.7000 7.5000 83.8000 ;
	    RECT 8.5000 83.7000 8.9000 83.8000 ;
	    RECT 5.4000 83.1000 5.8000 83.5000 ;
	    RECT 7.1000 83.4000 8.9000 83.7000 ;
	    RECT 7.5000 83.1000 7.8000 83.4000 ;
	    RECT 10.2000 83.1000 10.6000 83.5000 ;
	    RECT 5.1000 81.1000 5.7000 83.1000 ;
	    RECT 7.4000 81.1000 7.8000 83.1000 ;
	    RECT 9.6000 82.8000 10.6000 83.1000 ;
	    RECT 9.6000 81.1000 10.0000 82.8000 ;
	    RECT 11.8000 81.1000 12.2000 85.3000 ;
	    RECT 14.6000 85.1000 14.9000 85.8000 ;
	    RECT 15.3000 85.7000 15.7000 85.8000 ;
	    RECT 15.3000 85.4000 17.0000 85.7000 ;
	    RECT 16.7000 85.1000 17.0000 85.4000 ;
	    RECT 19.7000 85.1000 20.0000 86.8000 ;
	    RECT 22.4000 86.5000 22.7000 87.3000 ;
	    RECT 23.2000 87.2000 23.5000 87.9000 ;
	    RECT 24.6000 87.8000 25.0000 88.6000 ;
	    RECT 23.0000 86.8000 23.5000 87.2000 ;
	    RECT 22.4000 86.1000 22.9000 86.5000 ;
	    RECT 20.6000 85.1000 21.0000 85.2000 ;
	    RECT 22.4000 85.1000 22.7000 86.1000 ;
	    RECT 23.2000 85.1000 23.5000 86.8000 ;
	    RECT 12.6000 84.8000 13.8000 85.1000 ;
	    RECT 14.6000 84.8000 15.6000 85.1000 ;
	    RECT 12.6000 81.1000 13.0000 84.8000 ;
	    RECT 13.4000 84.7000 13.8000 84.8000 ;
	    RECT 14.8000 81.1000 15.6000 84.8000 ;
	    RECT 16.7000 84.8000 17.8000 85.1000 ;
	    RECT 16.7000 84.7000 17.1000 84.8000 ;
	    RECT 17.4000 81.1000 17.8000 84.8000 ;
	    RECT 19.5000 84.8000 20.0000 85.1000 ;
	    RECT 20.3000 84.8000 21.0000 85.1000 ;
	    RECT 21.4000 84.8000 22.7000 85.1000 ;
	    RECT 19.5000 82.2000 19.9000 84.8000 ;
	    RECT 20.3000 84.2000 20.6000 84.8000 ;
	    RECT 20.2000 83.8000 20.6000 84.2000 ;
	    RECT 19.0000 81.8000 19.9000 82.2000 ;
	    RECT 19.5000 81.1000 19.9000 81.8000 ;
	    RECT 21.4000 81.1000 21.8000 84.8000 ;
	    RECT 23.0000 84.6000 23.5000 85.1000 ;
	    RECT 25.4000 86.1000 25.8000 89.9000 ;
	    RECT 27.0000 88.8000 27.4000 89.9000 ;
	    RECT 27.0000 87.2000 27.3000 88.8000 ;
	    RECT 27.8000 87.8000 28.2000 88.6000 ;
	    RECT 28.6000 87.9000 29.0000 89.9000 ;
	    RECT 30.8000 88.1000 31.6000 89.9000 ;
	    RECT 28.6000 87.6000 29.8000 87.9000 ;
	    RECT 29.4000 87.5000 29.8000 87.6000 ;
	    RECT 30.1000 87.4000 30.5000 87.8000 ;
	    RECT 30.1000 87.2000 30.4000 87.4000 ;
	    RECT 27.0000 86.8000 27.4000 87.2000 ;
	    RECT 28.6000 86.8000 29.4000 87.2000 ;
	    RECT 30.0000 86.8000 30.4000 87.2000 ;
	    RECT 26.2000 86.1000 26.6000 86.2000 ;
	    RECT 25.4000 85.8000 26.6000 86.1000 ;
	    RECT 23.0000 81.1000 23.4000 84.6000 ;
	    RECT 25.4000 81.1000 25.8000 85.8000 ;
	    RECT 26.2000 85.4000 26.6000 85.8000 ;
	    RECT 27.0000 85.1000 27.3000 86.8000 ;
	    RECT 30.8000 86.4000 31.1000 88.1000 ;
	    RECT 33.4000 87.9000 33.8000 89.9000 ;
	    RECT 31.4000 87.7000 32.2000 87.8000 ;
	    RECT 31.4000 87.4000 32.4000 87.7000 ;
	    RECT 32.7000 87.6000 33.8000 87.9000 ;
	    RECT 32.7000 87.5000 33.1000 87.6000 ;
	    RECT 34.2000 87.5000 34.6000 89.9000 ;
	    RECT 36.4000 89.2000 36.8000 89.9000 ;
	    RECT 35.8000 88.9000 36.8000 89.2000 ;
	    RECT 38.6000 88.9000 39.0000 89.9000 ;
	    RECT 40.7000 89.2000 41.3000 89.9000 ;
	    RECT 40.6000 88.9000 41.3000 89.2000 ;
	    RECT 35.8000 88.5000 36.2000 88.9000 ;
	    RECT 38.6000 88.6000 38.9000 88.9000 ;
	    RECT 36.6000 88.2000 37.0000 88.6000 ;
	    RECT 37.5000 88.3000 38.9000 88.6000 ;
	    RECT 40.6000 88.5000 41.0000 88.9000 ;
	    RECT 37.5000 88.2000 37.9000 88.3000 ;
	    RECT 32.1000 87.2000 32.4000 87.4000 ;
	    RECT 31.4000 86.7000 31.8000 87.1000 ;
	    RECT 32.1000 86.9000 33.8000 87.2000 ;
	    RECT 33.0000 86.8000 33.8000 86.9000 ;
	    RECT 34.6000 87.1000 35.4000 87.2000 ;
	    RECT 36.7000 87.1000 37.0000 88.2000 ;
	    RECT 41.5000 87.7000 41.9000 87.8000 ;
	    RECT 43.0000 87.7000 43.4000 89.9000 ;
	    RECT 41.5000 87.4000 43.4000 87.7000 ;
	    RECT 39.5000 87.1000 39.9000 87.2000 ;
	    RECT 34.6000 86.8000 40.1000 87.1000 ;
	    RECT 36.1000 86.7000 36.5000 86.8000 ;
	    RECT 30.6000 86.2000 31.1000 86.4000 ;
	    RECT 30.2000 86.1000 31.1000 86.2000 ;
	    RECT 31.5000 86.4000 31.8000 86.7000 ;
	    RECT 31.5000 86.1000 32.8000 86.4000 ;
	    RECT 30.2000 85.8000 30.9000 86.1000 ;
	    RECT 32.4000 86.0000 32.8000 86.1000 ;
	    RECT 35.3000 86.2000 35.7000 86.3000 ;
	    RECT 35.3000 85.9000 37.8000 86.2000 ;
	    RECT 37.4000 85.8000 37.8000 85.9000 ;
	    RECT 30.6000 85.1000 30.9000 85.8000 ;
	    RECT 31.3000 85.7000 31.7000 85.8000 ;
	    RECT 31.3000 85.4000 33.0000 85.7000 ;
	    RECT 32.7000 85.1000 33.0000 85.4000 ;
	    RECT 34.2000 85.5000 37.0000 85.6000 ;
	    RECT 34.2000 85.4000 37.1000 85.5000 ;
	    RECT 34.2000 85.3000 39.1000 85.4000 ;
	    RECT 26.5000 84.7000 27.4000 85.1000 ;
	    RECT 28.6000 84.8000 29.8000 85.1000 ;
	    RECT 30.6000 84.8000 31.6000 85.1000 ;
	    RECT 26.5000 81.1000 26.9000 84.7000 ;
	    RECT 28.6000 81.1000 29.0000 84.8000 ;
	    RECT 29.4000 84.7000 29.8000 84.8000 ;
	    RECT 30.8000 84.2000 31.6000 84.8000 ;
	    RECT 32.7000 84.8000 33.8000 85.1000 ;
	    RECT 32.7000 84.7000 33.1000 84.8000 ;
	    RECT 30.2000 83.8000 31.6000 84.2000 ;
	    RECT 30.8000 81.1000 31.6000 83.8000 ;
	    RECT 33.4000 81.1000 33.8000 84.8000 ;
	    RECT 34.2000 81.1000 34.6000 85.3000 ;
	    RECT 36.7000 85.1000 39.1000 85.3000 ;
	    RECT 35.8000 84.5000 38.5000 84.8000 ;
	    RECT 35.8000 84.4000 36.2000 84.5000 ;
	    RECT 38.1000 84.4000 38.5000 84.5000 ;
	    RECT 38.8000 84.5000 39.1000 85.1000 ;
	    RECT 39.8000 85.2000 40.1000 86.8000 ;
	    RECT 40.6000 86.4000 41.0000 86.5000 ;
	    RECT 40.6000 86.1000 42.5000 86.4000 ;
	    RECT 42.1000 86.0000 42.5000 86.1000 ;
	    RECT 41.3000 85.7000 41.7000 85.8000 ;
	    RECT 43.0000 85.7000 43.4000 87.4000 ;
	    RECT 44.4000 87.1000 44.8000 89.9000 ;
	    RECT 48.6000 87.9000 49.0000 89.9000 ;
	    RECT 49.4000 88.0000 49.8000 89.9000 ;
	    RECT 51.0000 88.0000 51.4000 89.9000 ;
	    RECT 49.4000 87.9000 51.4000 88.0000 ;
	    RECT 51.8000 87.9000 52.2000 89.9000 ;
	    RECT 52.6000 88.0000 53.0000 89.9000 ;
	    RECT 54.2000 88.0000 54.6000 89.9000 ;
	    RECT 52.6000 87.9000 54.6000 88.0000 ;
	    RECT 48.7000 87.2000 49.0000 87.9000 ;
	    RECT 49.5000 87.7000 51.3000 87.9000 ;
	    RECT 50.6000 87.2000 51.0000 87.4000 ;
	    RECT 51.9000 87.2000 52.2000 87.9000 ;
	    RECT 52.7000 87.7000 54.5000 87.9000 ;
	    RECT 53.8000 87.2000 54.2000 87.4000 ;
	    RECT 41.3000 85.4000 43.4000 85.7000 ;
	    RECT 39.8000 84.9000 41.0000 85.2000 ;
	    RECT 39.5000 84.5000 39.9000 84.6000 ;
	    RECT 38.8000 84.2000 39.9000 84.5000 ;
	    RECT 40.7000 84.4000 41.0000 84.9000 ;
	    RECT 40.7000 84.0000 41.4000 84.4000 ;
	    RECT 37.5000 83.7000 37.9000 83.8000 ;
	    RECT 38.9000 83.7000 39.3000 83.8000 ;
	    RECT 35.8000 83.1000 36.2000 83.5000 ;
	    RECT 37.5000 83.4000 39.3000 83.7000 ;
	    RECT 38.6000 83.1000 38.9000 83.4000 ;
	    RECT 40.6000 83.1000 41.0000 83.5000 ;
	    RECT 35.8000 82.8000 36.8000 83.1000 ;
	    RECT 36.4000 81.1000 36.8000 82.8000 ;
	    RECT 38.6000 81.1000 39.0000 83.1000 ;
	    RECT 40.7000 81.1000 41.3000 83.1000 ;
	    RECT 43.0000 81.1000 43.4000 85.4000 ;
	    RECT 43.9000 86.9000 44.8000 87.1000 ;
	    RECT 47.8000 87.1000 48.2000 87.2000 ;
	    RECT 48.6000 87.1000 49.9000 87.2000 ;
	    RECT 43.9000 86.8000 44.7000 86.9000 ;
	    RECT 47.8000 86.8000 49.9000 87.1000 ;
	    RECT 50.6000 86.9000 51.4000 87.2000 ;
	    RECT 51.0000 86.8000 51.4000 86.9000 ;
	    RECT 51.8000 86.8000 53.1000 87.2000 ;
	    RECT 53.8000 86.9000 54.6000 87.2000 ;
	    RECT 54.2000 86.8000 54.6000 86.9000 ;
	    RECT 43.9000 85.2000 44.2000 86.8000 ;
	    RECT 45.0000 85.8000 45.8000 86.2000 ;
	    RECT 43.8000 84.8000 44.2000 85.2000 ;
	    RECT 46.2000 84.8000 46.6000 85.6000 ;
	    RECT 47.8000 85.1000 48.2000 85.2000 ;
	    RECT 48.6000 85.1000 49.0000 85.2000 ;
	    RECT 49.6000 85.1000 49.9000 86.8000 ;
	    RECT 50.2000 86.1000 50.6000 86.6000 ;
	    RECT 51.0000 86.1000 51.4000 86.2000 ;
	    RECT 50.2000 85.8000 51.4000 86.1000 ;
	    RECT 51.8000 85.1000 52.2000 85.2000 ;
	    RECT 52.8000 85.1000 53.1000 86.8000 ;
	    RECT 53.4000 85.8000 53.8000 86.6000 ;
	    RECT 54.2000 86.1000 54.6000 86.2000 ;
	    RECT 55.0000 86.1000 55.4000 89.9000 ;
	    RECT 56.6000 87.8000 57.0000 88.6000 ;
	    RECT 55.8000 87.1000 56.2000 87.6000 ;
	    RECT 56.6000 87.1000 57.0000 87.2000 ;
	    RECT 55.8000 86.8000 57.0000 87.1000 ;
	    RECT 54.2000 85.8000 55.4000 86.1000 ;
	    RECT 47.8000 84.8000 49.3000 85.1000 ;
	    RECT 49.6000 84.8000 50.1000 85.1000 ;
	    RECT 51.8000 84.8000 52.5000 85.1000 ;
	    RECT 52.8000 84.8000 53.3000 85.1000 ;
	    RECT 43.9000 83.5000 44.2000 84.8000 ;
	    RECT 44.6000 83.8000 45.0000 84.6000 ;
	    RECT 49.0000 84.2000 49.3000 84.8000 ;
	    RECT 49.0000 83.8000 49.4000 84.2000 ;
	    RECT 43.9000 83.2000 45.7000 83.5000 ;
	    RECT 43.9000 83.1000 44.2000 83.2000 ;
	    RECT 43.8000 81.1000 44.2000 83.1000 ;
	    RECT 45.4000 81.1000 45.8000 83.2000 ;
	    RECT 49.7000 81.1000 50.1000 84.8000 ;
	    RECT 52.2000 84.2000 52.5000 84.8000 ;
	    RECT 52.2000 83.8000 52.6000 84.2000 ;
	    RECT 52.9000 81.1000 53.3000 84.8000 ;
	    RECT 55.0000 81.1000 55.4000 85.8000 ;
	    RECT 57.4000 81.1000 57.8000 89.9000 ;
	    RECT 58.8000 89.2000 59.2000 89.9000 ;
	    RECT 61.7000 89.2000 62.1000 89.9000 ;
	    RECT 58.2000 88.8000 59.2000 89.2000 ;
	    RECT 61.4000 88.8000 62.1000 89.2000 ;
	    RECT 58.8000 87.1000 59.2000 88.8000 ;
	    RECT 61.7000 88.4000 62.1000 88.8000 ;
	    RECT 58.3000 86.9000 59.2000 87.1000 ;
	    RECT 61.4000 87.9000 62.1000 88.4000 ;
	    RECT 63.8000 87.9000 64.2000 89.9000 ;
	    RECT 58.3000 86.8000 59.1000 86.9000 ;
	    RECT 58.3000 85.2000 58.6000 86.8000 ;
	    RECT 61.4000 86.2000 61.7000 87.9000 ;
	    RECT 63.8000 87.8000 64.1000 87.9000 ;
	    RECT 63.2000 87.6000 64.1000 87.8000 ;
	    RECT 62.0000 87.5000 64.1000 87.6000 ;
	    RECT 62.0000 87.3000 63.5000 87.5000 ;
	    RECT 62.0000 87.2000 62.4000 87.3000 ;
	    RECT 59.0000 85.8000 60.2000 86.2000 ;
	    RECT 61.4000 85.8000 61.8000 86.2000 ;
	    RECT 58.2000 84.8000 58.6000 85.2000 ;
	    RECT 60.6000 84.8000 61.0000 85.6000 ;
	    RECT 61.4000 85.1000 61.7000 85.8000 ;
	    RECT 62.1000 85.5000 62.4000 87.2000 ;
	    RECT 62.8000 86.9000 63.2000 87.0000 ;
	    RECT 62.8000 86.6000 63.3000 86.9000 ;
	    RECT 63.0000 86.2000 63.3000 86.6000 ;
	    RECT 63.8000 86.4000 64.2000 87.2000 ;
	    RECT 63.0000 85.8000 63.4000 86.2000 ;
	    RECT 62.1000 85.2000 63.3000 85.5000 ;
	    RECT 58.3000 83.5000 58.6000 84.8000 ;
	    RECT 59.0000 83.8000 59.4000 84.6000 ;
	    RECT 58.3000 83.2000 60.1000 83.5000 ;
	    RECT 58.3000 83.1000 58.6000 83.2000 ;
	    RECT 58.2000 81.1000 58.6000 83.1000 ;
	    RECT 59.8000 83.1000 60.1000 83.2000 ;
	    RECT 59.8000 81.1000 60.2000 83.1000 ;
	    RECT 61.4000 81.1000 61.8000 85.1000 ;
	    RECT 63.0000 83.1000 63.3000 85.2000 ;
	    RECT 63.8000 85.1000 64.2000 85.2000 ;
	    RECT 64.6000 85.1000 65.0000 89.9000 ;
	    RECT 65.4000 87.8000 65.8000 88.6000 ;
	    RECT 66.2000 88.0000 66.6000 89.9000 ;
	    RECT 67.8000 88.0000 68.2000 89.9000 ;
	    RECT 66.2000 87.9000 68.2000 88.0000 ;
	    RECT 68.6000 87.9000 69.0000 89.9000 ;
	    RECT 70.2000 88.2000 70.6000 89.9000 ;
	    RECT 70.1000 87.9000 70.6000 88.2000 ;
	    RECT 66.3000 87.7000 68.1000 87.9000 ;
	    RECT 66.6000 87.2000 67.0000 87.4000 ;
	    RECT 68.6000 87.2000 68.9000 87.9000 ;
	    RECT 70.1000 87.2000 70.4000 87.9000 ;
	    RECT 71.8000 87.6000 72.2000 89.9000 ;
	    RECT 72.6000 87.9000 73.0000 89.9000 ;
	    RECT 74.8000 89.2000 75.6000 89.9000 ;
	    RECT 74.8000 88.8000 76.2000 89.2000 ;
	    RECT 74.8000 88.1000 75.6000 88.8000 ;
	    RECT 72.6000 87.6000 73.7000 87.9000 ;
	    RECT 74.2000 87.7000 75.0000 87.8000 ;
	    RECT 70.9000 87.3000 72.2000 87.6000 ;
	    RECT 73.3000 87.5000 73.7000 87.6000 ;
	    RECT 74.0000 87.4000 75.0000 87.7000 ;
	    RECT 66.2000 86.9000 67.0000 87.2000 ;
	    RECT 67.7000 87.1000 69.0000 87.2000 ;
	    RECT 66.2000 86.8000 66.6000 86.9000 ;
	    RECT 67.7000 86.8000 69.7000 87.1000 ;
	    RECT 65.4000 86.1000 65.8000 86.2000 ;
	    RECT 67.0000 86.1000 67.4000 86.6000 ;
	    RECT 65.4000 85.8000 67.4000 86.1000 ;
	    RECT 67.7000 85.1000 68.0000 86.8000 ;
	    RECT 69.4000 86.2000 69.7000 86.8000 ;
	    RECT 70.1000 86.8000 70.6000 87.2000 ;
	    RECT 69.4000 85.8000 69.8000 86.2000 ;
	    RECT 68.6000 85.1000 69.0000 85.2000 ;
	    RECT 63.8000 84.8000 65.0000 85.1000 ;
	    RECT 63.0000 81.1000 63.4000 83.1000 ;
	    RECT 64.6000 81.1000 65.0000 84.8000 ;
	    RECT 67.5000 84.8000 68.0000 85.1000 ;
	    RECT 68.3000 84.8000 69.0000 85.1000 ;
	    RECT 70.1000 85.1000 70.4000 86.8000 ;
	    RECT 70.9000 86.5000 71.2000 87.3000 ;
	    RECT 74.0000 87.2000 74.3000 87.4000 ;
	    RECT 72.6000 86.9000 74.3000 87.2000 ;
	    RECT 72.6000 86.8000 73.4000 86.9000 ;
	    RECT 74.6000 86.7000 75.0000 87.1000 ;
	    RECT 70.7000 86.1000 71.2000 86.5000 ;
	    RECT 70.9000 85.1000 71.2000 86.1000 ;
	    RECT 71.7000 86.2000 72.1000 86.6000 ;
	    RECT 74.6000 86.4000 74.9000 86.7000 ;
	    RECT 71.7000 85.8000 72.2000 86.2000 ;
	    RECT 73.6000 86.1000 74.9000 86.4000 ;
	    RECT 75.3000 86.4000 75.6000 88.1000 ;
	    RECT 77.4000 87.9000 77.8000 89.9000 ;
	    RECT 75.9000 87.4000 76.3000 87.8000 ;
	    RECT 76.6000 87.6000 77.8000 87.9000 ;
	    RECT 78.2000 87.7000 78.6000 89.9000 ;
	    RECT 80.3000 89.2000 80.9000 89.9000 ;
	    RECT 80.3000 88.9000 81.0000 89.2000 ;
	    RECT 82.6000 88.9000 83.0000 89.9000 ;
	    RECT 84.8000 89.2000 85.2000 89.9000 ;
	    RECT 84.8000 88.9000 85.8000 89.2000 ;
	    RECT 80.6000 88.5000 81.0000 88.9000 ;
	    RECT 82.7000 88.6000 83.0000 88.9000 ;
	    RECT 82.7000 88.3000 84.1000 88.6000 ;
	    RECT 83.7000 88.2000 84.1000 88.3000 ;
	    RECT 84.6000 88.2000 85.0000 88.6000 ;
	    RECT 85.4000 88.5000 85.8000 88.9000 ;
	    RECT 79.7000 87.7000 80.1000 87.8000 ;
	    RECT 76.6000 87.5000 77.0000 87.6000 ;
	    RECT 76.0000 87.2000 76.3000 87.4000 ;
	    RECT 78.2000 87.4000 80.1000 87.7000 ;
	    RECT 76.0000 86.8000 76.4000 87.2000 ;
	    RECT 77.0000 86.8000 77.8000 87.2000 ;
	    RECT 75.3000 86.2000 75.8000 86.4000 ;
	    RECT 75.3000 86.1000 76.2000 86.2000 ;
	    RECT 73.6000 86.0000 74.0000 86.1000 ;
	    RECT 75.5000 85.8000 76.2000 86.1000 ;
	    RECT 74.7000 85.7000 75.1000 85.8000 ;
	    RECT 73.4000 85.4000 75.1000 85.7000 ;
	    RECT 73.4000 85.1000 73.7000 85.4000 ;
	    RECT 75.5000 85.1000 75.8000 85.8000 ;
	    RECT 78.2000 85.7000 78.6000 87.4000 ;
	    RECT 81.7000 87.1000 82.1000 87.2000 ;
	    RECT 84.6000 87.1000 84.9000 88.2000 ;
	    RECT 87.0000 87.5000 87.4000 89.9000 ;
	    RECT 87.8000 87.6000 88.2000 89.9000 ;
	    RECT 89.4000 88.2000 89.8000 89.9000 ;
	    RECT 89.4000 87.9000 89.9000 88.2000 ;
	    RECT 87.8000 87.3000 89.1000 87.6000 ;
	    RECT 86.2000 87.1000 87.0000 87.2000 ;
	    RECT 81.5000 86.8000 87.0000 87.1000 ;
	    RECT 80.6000 86.4000 81.0000 86.5000 ;
	    RECT 79.1000 86.1000 81.0000 86.4000 ;
	    RECT 79.1000 86.0000 79.5000 86.1000 ;
	    RECT 79.9000 85.7000 80.3000 85.8000 ;
	    RECT 78.2000 85.4000 80.3000 85.7000 ;
	    RECT 67.5000 81.1000 67.9000 84.8000 ;
	    RECT 68.3000 84.2000 68.6000 84.8000 ;
	    RECT 70.1000 84.6000 70.6000 85.1000 ;
	    RECT 70.9000 84.8000 72.2000 85.1000 ;
	    RECT 68.2000 83.8000 68.6000 84.2000 ;
	    RECT 70.2000 81.1000 70.6000 84.6000 ;
	    RECT 71.8000 81.1000 72.2000 84.8000 ;
	    RECT 72.6000 84.8000 73.7000 85.1000 ;
	    RECT 72.6000 81.1000 73.0000 84.8000 ;
	    RECT 73.3000 84.7000 73.7000 84.8000 ;
	    RECT 74.8000 84.8000 75.8000 85.1000 ;
	    RECT 76.6000 84.8000 77.8000 85.1000 ;
	    RECT 74.8000 81.1000 75.6000 84.8000 ;
	    RECT 76.6000 84.7000 77.0000 84.8000 ;
	    RECT 77.4000 81.1000 77.8000 84.8000 ;
	    RECT 78.2000 81.1000 78.6000 85.4000 ;
	    RECT 81.5000 85.2000 81.8000 86.8000 ;
	    RECT 85.1000 86.7000 85.5000 86.8000 ;
	    RECT 85.9000 86.2000 86.3000 86.3000 ;
	    RECT 87.9000 86.2000 88.3000 86.6000 ;
	    RECT 83.8000 85.9000 86.3000 86.2000 ;
	    RECT 83.8000 85.8000 84.2000 85.9000 ;
	    RECT 87.8000 85.8000 88.3000 86.2000 ;
	    RECT 88.8000 86.5000 89.1000 87.3000 ;
	    RECT 89.6000 87.2000 89.9000 87.9000 ;
	    RECT 91.0000 87.6000 91.4000 89.9000 ;
	    RECT 91.0000 87.3000 92.1000 87.6000 ;
	    RECT 89.4000 87.1000 89.9000 87.2000 ;
	    RECT 89.4000 86.8000 90.5000 87.1000 ;
	    RECT 88.8000 86.1000 89.3000 86.5000 ;
	    RECT 84.6000 85.5000 87.4000 85.6000 ;
	    RECT 84.5000 85.4000 87.4000 85.5000 ;
	    RECT 80.6000 84.9000 81.8000 85.2000 ;
	    RECT 82.5000 85.3000 87.4000 85.4000 ;
	    RECT 82.5000 85.1000 84.9000 85.3000 ;
	    RECT 80.6000 84.4000 80.9000 84.9000 ;
	    RECT 80.2000 84.2000 80.9000 84.4000 ;
	    RECT 81.7000 84.5000 82.1000 84.6000 ;
	    RECT 82.5000 84.5000 82.8000 85.1000 ;
	    RECT 81.7000 84.2000 82.8000 84.5000 ;
	    RECT 83.1000 84.5000 85.8000 84.8000 ;
	    RECT 83.1000 84.4000 83.5000 84.5000 ;
	    RECT 85.4000 84.4000 85.8000 84.5000 ;
	    RECT 79.8000 84.0000 80.9000 84.2000 ;
	    RECT 79.8000 83.8000 80.5000 84.0000 ;
	    RECT 82.3000 83.7000 82.7000 83.8000 ;
	    RECT 83.7000 83.7000 84.1000 83.8000 ;
	    RECT 80.6000 83.1000 81.0000 83.5000 ;
	    RECT 82.3000 83.4000 84.1000 83.7000 ;
	    RECT 82.7000 83.1000 83.0000 83.4000 ;
	    RECT 85.4000 83.1000 85.8000 83.5000 ;
	    RECT 80.3000 81.1000 80.9000 83.1000 ;
	    RECT 82.6000 81.1000 83.0000 83.1000 ;
	    RECT 84.8000 82.8000 85.8000 83.1000 ;
	    RECT 84.8000 81.1000 85.2000 82.8000 ;
	    RECT 87.0000 81.1000 87.4000 85.3000 ;
	    RECT 88.8000 85.1000 89.1000 86.1000 ;
	    RECT 89.6000 85.1000 89.9000 86.8000 ;
	    RECT 90.2000 86.1000 90.5000 86.8000 ;
	    RECT 91.0000 86.1000 91.4000 86.6000 ;
	    RECT 90.2000 85.8000 91.4000 86.1000 ;
	    RECT 91.8000 85.8000 92.1000 87.3000 ;
	    RECT 92.6000 86.2000 93.0000 89.9000 ;
	    RECT 93.4000 87.6000 93.8000 89.9000 ;
	    RECT 95.0000 88.2000 95.4000 89.9000 ;
	    RECT 95.0000 87.9000 95.5000 88.2000 ;
	    RECT 96.6000 87.9000 97.0000 89.9000 ;
	    RECT 97.4000 88.0000 97.8000 89.9000 ;
	    RECT 99.0000 88.0000 99.4000 89.9000 ;
	    RECT 97.4000 87.9000 99.4000 88.0000 ;
	    RECT 93.4000 87.3000 94.7000 87.6000 ;
	    RECT 91.8000 85.4000 92.4000 85.8000 ;
	    RECT 91.8000 85.1000 92.1000 85.4000 ;
	    RECT 92.7000 85.1000 93.0000 86.2000 ;
	    RECT 94.4000 86.5000 94.7000 87.3000 ;
	    RECT 95.2000 87.2000 95.5000 87.9000 ;
	    RECT 96.7000 87.2000 97.0000 87.9000 ;
	    RECT 97.5000 87.7000 99.3000 87.9000 ;
	    RECT 101.4000 87.6000 101.8000 89.9000 ;
	    RECT 103.0000 88.2000 103.4000 89.9000 ;
	    RECT 103.0000 87.9000 103.5000 88.2000 ;
	    RECT 98.6000 87.2000 99.0000 87.4000 ;
	    RECT 101.4000 87.3000 102.7000 87.6000 ;
	    RECT 95.0000 87.1000 95.5000 87.2000 ;
	    RECT 95.8000 87.1000 96.2000 87.2000 ;
	    RECT 95.0000 86.8000 96.2000 87.1000 ;
	    RECT 96.6000 86.8000 97.9000 87.2000 ;
	    RECT 98.6000 86.9000 99.4000 87.2000 ;
	    RECT 99.0000 86.8000 99.4000 86.9000 ;
	    RECT 94.4000 86.1000 94.9000 86.5000 ;
	    RECT 94.4000 85.1000 94.7000 86.1000 ;
	    RECT 95.2000 85.1000 95.5000 86.8000 ;
	    RECT 87.8000 84.8000 89.1000 85.1000 ;
	    RECT 87.8000 81.1000 88.2000 84.8000 ;
	    RECT 89.4000 84.6000 89.9000 85.1000 ;
	    RECT 91.0000 84.8000 92.1000 85.1000 ;
	    RECT 89.4000 81.1000 89.8000 84.6000 ;
	    RECT 91.0000 81.1000 91.4000 84.8000 ;
	    RECT 92.6000 81.1000 93.0000 85.1000 ;
	    RECT 93.4000 84.8000 94.7000 85.1000 ;
	    RECT 93.4000 81.1000 93.8000 84.8000 ;
	    RECT 95.0000 84.6000 95.5000 85.1000 ;
	    RECT 96.6000 85.1000 97.0000 85.2000 ;
	    RECT 97.6000 85.1000 97.9000 86.8000 ;
	    RECT 98.2000 85.8000 98.6000 86.6000 ;
	    RECT 102.4000 86.5000 102.7000 87.3000 ;
	    RECT 103.2000 87.2000 103.5000 87.9000 ;
	    RECT 103.0000 86.8000 103.5000 87.2000 ;
	    RECT 103.8000 87.1000 104.2000 87.2000 ;
	    RECT 104.6000 87.1000 105.0000 87.6000 ;
	    RECT 103.8000 86.8000 105.0000 87.1000 ;
	    RECT 102.4000 86.1000 102.9000 86.5000 ;
	    RECT 102.4000 85.1000 102.7000 86.1000 ;
	    RECT 103.2000 85.1000 103.5000 86.8000 ;
	    RECT 96.6000 84.8000 97.3000 85.1000 ;
	    RECT 97.6000 84.8000 98.1000 85.1000 ;
	    RECT 95.0000 81.1000 95.4000 84.6000 ;
	    RECT 97.0000 84.2000 97.3000 84.8000 ;
	    RECT 97.0000 83.8000 97.4000 84.2000 ;
	    RECT 97.7000 81.1000 98.1000 84.8000 ;
	    RECT 101.4000 84.8000 102.7000 85.1000 ;
	    RECT 101.4000 81.1000 101.8000 84.8000 ;
	    RECT 103.0000 84.6000 103.5000 85.1000 ;
	    RECT 105.4000 86.1000 105.8000 89.9000 ;
	    RECT 107.0000 88.0000 107.4000 89.9000 ;
	    RECT 108.6000 88.0000 109.0000 89.9000 ;
	    RECT 107.0000 87.9000 109.0000 88.0000 ;
	    RECT 109.4000 87.9000 109.8000 89.9000 ;
	    RECT 110.2000 87.9000 110.6000 89.9000 ;
	    RECT 112.3000 88.4000 112.7000 89.9000 ;
	    RECT 113.4000 89.6000 115.4000 89.9000 ;
	    RECT 112.3000 87.9000 113.0000 88.4000 ;
	    RECT 113.4000 87.9000 113.8000 89.6000 ;
	    RECT 114.2000 87.9000 114.6000 89.3000 ;
	    RECT 115.0000 88.0000 115.4000 89.6000 ;
	    RECT 116.6000 88.0000 117.0000 89.9000 ;
	    RECT 115.0000 87.9000 117.0000 88.0000 ;
	    RECT 107.1000 87.7000 108.9000 87.9000 ;
	    RECT 107.4000 87.2000 107.8000 87.4000 ;
	    RECT 109.4000 87.2000 109.7000 87.9000 ;
	    RECT 110.3000 87.8000 110.6000 87.9000 ;
	    RECT 110.3000 87.6000 111.2000 87.8000 ;
	    RECT 110.3000 87.5000 112.4000 87.6000 ;
	    RECT 110.9000 87.3000 112.4000 87.5000 ;
	    RECT 112.0000 87.2000 112.4000 87.3000 ;
	    RECT 107.0000 86.9000 107.8000 87.2000 ;
	    RECT 107.0000 86.8000 107.4000 86.9000 ;
	    RECT 108.5000 86.8000 109.8000 87.2000 ;
	    RECT 107.8000 86.1000 108.2000 86.6000 ;
	    RECT 105.4000 85.8000 108.2000 86.1000 ;
	    RECT 103.0000 81.1000 103.4000 84.6000 ;
	    RECT 105.4000 81.1000 105.8000 85.8000 ;
	    RECT 108.5000 85.2000 108.8000 86.8000 ;
	    RECT 110.2000 86.4000 110.6000 87.2000 ;
	    RECT 111.2000 86.9000 111.6000 87.0000 ;
	    RECT 111.1000 86.6000 111.6000 86.9000 ;
	    RECT 111.1000 86.2000 111.4000 86.6000 ;
	    RECT 111.0000 85.8000 111.4000 86.2000 ;
	    RECT 112.0000 85.5000 112.3000 87.2000 ;
	    RECT 112.7000 86.2000 113.0000 87.9000 ;
	    RECT 114.2000 87.2000 114.5000 87.9000 ;
	    RECT 115.1000 87.7000 116.9000 87.9000 ;
	    RECT 116.2000 87.2000 116.6000 87.4000 ;
	    RECT 112.6000 86.1000 113.0000 86.2000 ;
	    RECT 113.4000 86.1000 113.8000 87.2000 ;
	    RECT 114.2000 86.9000 115.4000 87.2000 ;
	    RECT 116.2000 86.9000 117.0000 87.2000 ;
	    RECT 118.0000 87.1000 118.4000 89.9000 ;
	    RECT 115.0000 86.8000 115.4000 86.9000 ;
	    RECT 116.6000 86.8000 117.0000 86.9000 ;
	    RECT 117.5000 86.9000 118.4000 87.1000 ;
	    RECT 117.5000 86.8000 118.3000 86.9000 ;
	    RECT 120.6000 86.8000 121.0000 87.6000 ;
	    RECT 112.6000 85.8000 113.8000 86.1000 ;
	    RECT 114.2000 85.8000 114.6000 86.6000 ;
	    RECT 111.1000 85.2000 112.3000 85.5000 ;
	    RECT 108.4000 85.1000 108.8000 85.2000 ;
	    RECT 109.4000 85.1000 109.8000 85.2000 ;
	    RECT 108.3000 84.8000 108.8000 85.1000 ;
	    RECT 109.1000 84.8000 109.8000 85.1000 ;
	    RECT 108.3000 81.1000 108.7000 84.8000 ;
	    RECT 109.1000 84.2000 109.4000 84.8000 ;
	    RECT 109.0000 83.8000 109.4000 84.2000 ;
	    RECT 111.1000 83.1000 111.4000 85.2000 ;
	    RECT 112.7000 85.1000 113.0000 85.8000 ;
	    RECT 115.1000 85.1000 115.4000 86.8000 ;
	    RECT 115.8000 85.8000 116.2000 86.6000 ;
	    RECT 117.5000 85.2000 117.8000 86.8000 ;
	    RECT 118.6000 85.8000 119.4000 86.2000 ;
	    RECT 111.0000 81.1000 111.4000 83.1000 ;
	    RECT 112.6000 81.1000 113.0000 85.1000 ;
	    RECT 114.7000 81.1000 115.7000 85.1000 ;
	    RECT 117.4000 84.8000 117.8000 85.2000 ;
	    RECT 119.8000 84.8000 120.2000 85.6000 ;
	    RECT 117.5000 83.5000 117.8000 84.8000 ;
	    RECT 118.2000 83.8000 118.6000 84.6000 ;
	    RECT 117.5000 83.2000 119.3000 83.5000 ;
	    RECT 117.5000 83.1000 117.8000 83.2000 ;
	    RECT 117.4000 81.1000 117.8000 83.1000 ;
	    RECT 119.0000 83.1000 119.3000 83.2000 ;
	    RECT 119.0000 81.1000 119.4000 83.1000 ;
	    RECT 121.4000 81.1000 121.8000 89.9000 ;
	    RECT 123.0000 87.7000 123.4000 89.9000 ;
	    RECT 125.1000 89.2000 125.7000 89.9000 ;
	    RECT 125.1000 88.9000 125.8000 89.2000 ;
	    RECT 127.4000 88.9000 127.8000 89.9000 ;
	    RECT 129.6000 89.2000 130.0000 89.9000 ;
	    RECT 129.6000 88.9000 130.6000 89.2000 ;
	    RECT 125.4000 88.5000 125.8000 88.9000 ;
	    RECT 127.5000 88.6000 127.8000 88.9000 ;
	    RECT 127.5000 88.3000 128.9000 88.6000 ;
	    RECT 128.5000 88.2000 128.9000 88.3000 ;
	    RECT 129.4000 88.2000 129.8000 88.6000 ;
	    RECT 130.2000 88.5000 130.6000 88.9000 ;
	    RECT 124.5000 87.7000 124.9000 87.8000 ;
	    RECT 123.0000 87.4000 124.9000 87.7000 ;
	    RECT 123.0000 85.7000 123.4000 87.4000 ;
	    RECT 126.5000 87.1000 126.9000 87.2000 ;
	    RECT 129.4000 87.1000 129.7000 88.2000 ;
	    RECT 131.8000 87.5000 132.2000 89.9000 ;
	    RECT 132.6000 87.5000 133.0000 89.9000 ;
	    RECT 134.8000 89.2000 135.2000 89.9000 ;
	    RECT 134.2000 88.9000 135.2000 89.2000 ;
	    RECT 137.0000 88.9000 137.4000 89.9000 ;
	    RECT 139.1000 89.2000 139.7000 89.9000 ;
	    RECT 139.0000 88.9000 139.7000 89.2000 ;
	    RECT 134.2000 88.5000 134.6000 88.9000 ;
	    RECT 137.0000 88.6000 137.3000 88.9000 ;
	    RECT 135.0000 88.2000 135.4000 88.6000 ;
	    RECT 135.9000 88.3000 137.3000 88.6000 ;
	    RECT 139.0000 88.5000 139.4000 88.9000 ;
	    RECT 135.9000 88.2000 136.3000 88.3000 ;
	    RECT 131.0000 87.1000 131.8000 87.2000 ;
	    RECT 133.0000 87.1000 133.8000 87.2000 ;
	    RECT 135.1000 87.1000 135.4000 88.2000 ;
	    RECT 139.9000 87.7000 140.3000 87.8000 ;
	    RECT 141.4000 87.7000 141.8000 89.9000 ;
	    RECT 143.0000 88.2000 143.4000 89.9000 ;
	    RECT 139.9000 87.4000 141.8000 87.7000 ;
	    RECT 137.9000 87.1000 138.3000 87.2000 ;
	    RECT 126.3000 86.8000 138.5000 87.1000 ;
	    RECT 125.4000 86.4000 125.8000 86.5000 ;
	    RECT 123.9000 86.1000 125.8000 86.4000 ;
	    RECT 123.9000 86.0000 124.3000 86.1000 ;
	    RECT 124.7000 85.7000 125.1000 85.8000 ;
	    RECT 123.0000 85.4000 125.1000 85.7000 ;
	    RECT 123.0000 81.1000 123.4000 85.4000 ;
	    RECT 126.3000 85.2000 126.6000 86.8000 ;
	    RECT 129.9000 86.7000 130.3000 86.8000 ;
	    RECT 134.5000 86.7000 134.9000 86.8000 ;
	    RECT 129.4000 86.2000 129.8000 86.3000 ;
	    RECT 130.7000 86.2000 131.1000 86.3000 ;
	    RECT 128.6000 85.9000 131.1000 86.2000 ;
	    RECT 133.7000 86.2000 134.1000 86.3000 ;
	    RECT 135.0000 86.2000 135.4000 86.3000 ;
	    RECT 133.7000 85.9000 136.2000 86.2000 ;
	    RECT 128.6000 85.8000 129.0000 85.9000 ;
	    RECT 135.8000 85.8000 136.2000 85.9000 ;
	    RECT 129.4000 85.5000 132.2000 85.6000 ;
	    RECT 129.3000 85.4000 132.2000 85.5000 ;
	    RECT 125.4000 84.9000 126.6000 85.2000 ;
	    RECT 127.3000 85.3000 132.2000 85.4000 ;
	    RECT 127.3000 85.1000 129.7000 85.3000 ;
	    RECT 125.4000 84.4000 125.7000 84.9000 ;
	    RECT 125.0000 84.0000 125.7000 84.4000 ;
	    RECT 126.5000 84.5000 126.9000 84.6000 ;
	    RECT 127.3000 84.5000 127.6000 85.1000 ;
	    RECT 126.5000 84.2000 127.6000 84.5000 ;
	    RECT 127.9000 84.5000 130.6000 84.8000 ;
	    RECT 127.9000 84.4000 128.3000 84.5000 ;
	    RECT 130.2000 84.4000 130.6000 84.5000 ;
	    RECT 127.1000 83.7000 127.5000 83.8000 ;
	    RECT 128.5000 83.7000 128.9000 83.8000 ;
	    RECT 125.4000 83.1000 125.8000 83.5000 ;
	    RECT 127.1000 83.4000 128.9000 83.7000 ;
	    RECT 127.5000 83.1000 127.8000 83.4000 ;
	    RECT 130.2000 83.1000 130.6000 83.5000 ;
	    RECT 125.1000 81.1000 125.7000 83.1000 ;
	    RECT 127.4000 81.1000 127.8000 83.1000 ;
	    RECT 129.6000 82.8000 130.6000 83.1000 ;
	    RECT 129.6000 81.1000 130.0000 82.8000 ;
	    RECT 131.8000 81.1000 132.2000 85.3000 ;
	    RECT 132.6000 85.5000 135.4000 85.6000 ;
	    RECT 132.6000 85.4000 135.5000 85.5000 ;
	    RECT 132.6000 85.3000 137.5000 85.4000 ;
	    RECT 132.6000 81.1000 133.0000 85.3000 ;
	    RECT 135.1000 85.1000 137.5000 85.3000 ;
	    RECT 134.2000 84.5000 136.9000 84.8000 ;
	    RECT 134.2000 84.4000 134.6000 84.5000 ;
	    RECT 136.5000 84.4000 136.9000 84.5000 ;
	    RECT 137.2000 84.5000 137.5000 85.1000 ;
	    RECT 138.2000 85.2000 138.5000 86.8000 ;
	    RECT 139.0000 86.4000 139.4000 86.5000 ;
	    RECT 139.0000 86.1000 140.9000 86.4000 ;
	    RECT 140.5000 86.0000 140.9000 86.1000 ;
	    RECT 139.7000 85.7000 140.1000 85.8000 ;
	    RECT 141.4000 85.7000 141.8000 87.4000 ;
	    RECT 139.7000 85.4000 141.8000 85.7000 ;
	    RECT 138.2000 84.9000 139.4000 85.2000 ;
	    RECT 137.9000 84.5000 138.3000 84.6000 ;
	    RECT 137.2000 84.2000 138.3000 84.5000 ;
	    RECT 139.1000 84.4000 139.4000 84.9000 ;
	    RECT 139.1000 84.0000 139.8000 84.4000 ;
	    RECT 135.9000 83.7000 136.3000 83.8000 ;
	    RECT 137.3000 83.7000 137.7000 83.8000 ;
	    RECT 134.2000 83.1000 134.6000 83.5000 ;
	    RECT 135.9000 83.4000 137.7000 83.7000 ;
	    RECT 137.0000 83.1000 137.3000 83.4000 ;
	    RECT 139.0000 83.1000 139.4000 83.5000 ;
	    RECT 134.2000 82.8000 135.2000 83.1000 ;
	    RECT 134.8000 81.1000 135.2000 82.8000 ;
	    RECT 137.0000 81.1000 137.4000 83.1000 ;
	    RECT 139.1000 81.1000 139.7000 83.1000 ;
	    RECT 141.4000 81.1000 141.8000 85.4000 ;
	    RECT 142.9000 87.9000 143.4000 88.2000 ;
	    RECT 142.9000 87.2000 143.2000 87.9000 ;
	    RECT 144.6000 87.6000 145.0000 89.9000 ;
	    RECT 143.7000 87.3000 145.0000 87.6000 ;
	    RECT 145.4000 87.6000 145.8000 89.9000 ;
	    RECT 145.4000 87.3000 146.5000 87.6000 ;
	    RECT 142.9000 86.8000 143.4000 87.2000 ;
	    RECT 142.9000 85.1000 143.2000 86.8000 ;
	    RECT 143.7000 86.5000 144.0000 87.3000 ;
	    RECT 143.5000 86.1000 144.0000 86.5000 ;
	    RECT 143.7000 85.1000 144.0000 86.1000 ;
	    RECT 144.5000 86.2000 144.9000 86.6000 ;
	    RECT 144.5000 85.8000 145.0000 86.2000 ;
	    RECT 145.4000 85.8000 145.8000 86.6000 ;
	    RECT 146.2000 85.8000 146.5000 87.3000 ;
	    RECT 146.2000 85.4000 146.8000 85.8000 ;
	    RECT 146.2000 85.1000 146.5000 85.4000 ;
	    RECT 142.9000 84.6000 143.4000 85.1000 ;
	    RECT 143.7000 84.8000 145.0000 85.1000 ;
	    RECT 143.0000 81.1000 143.4000 84.6000 ;
	    RECT 144.6000 81.1000 145.0000 84.8000 ;
	    RECT 145.4000 84.8000 146.5000 85.1000 ;
	    RECT 145.4000 81.1000 145.8000 84.8000 ;
	    RECT 2.2000 76.2000 2.6000 79.9000 ;
	    RECT 3.1000 79.6000 4.9000 79.9000 ;
	    RECT 3.1000 79.5000 3.4000 79.6000 ;
	    RECT 3.0000 76.5000 3.4000 79.5000 ;
	    RECT 4.6000 79.5000 4.9000 79.6000 ;
	    RECT 5.4000 79.6000 7.4000 79.9000 ;
	    RECT 3.8000 76.5000 4.2000 79.3000 ;
	    RECT 4.6000 76.7000 5.0000 79.5000 ;
	    RECT 5.4000 77.0000 5.8000 79.6000 ;
	    RECT 6.2000 76.9000 6.6000 79.3000 ;
	    RECT 7.0000 76.9000 7.4000 79.6000 ;
	    RECT 6.2000 76.7000 6.5000 76.9000 ;
	    RECT 4.6000 76.5000 6.5000 76.7000 ;
	    RECT 3.9000 76.2000 4.2000 76.5000 ;
	    RECT 4.7000 76.4000 6.5000 76.5000 ;
	    RECT 7.1000 76.6000 7.4000 76.9000 ;
	    RECT 8.6000 76.9000 9.0000 79.9000 ;
	    RECT 10.2000 77.9000 10.6000 79.9000 ;
	    RECT 8.6000 76.6000 8.9000 76.9000 ;
	    RECT 7.1000 76.3000 8.9000 76.6000 ;
	    RECT 1.5000 75.9000 2.6000 76.2000 ;
	    RECT 3.8000 76.1000 4.2000 76.2000 ;
	    RECT 1.5000 75.6000 1.8000 75.9000 ;
	    RECT 3.8000 75.8000 5.5000 76.1000 ;
	    RECT 1.2000 75.2000 1.8000 75.6000 ;
	    RECT 1.5000 73.7000 1.8000 75.2000 ;
	    RECT 2.2000 75.1000 2.6000 75.2000 ;
	    RECT 3.8000 75.1000 4.2000 75.2000 ;
	    RECT 2.2000 74.8000 4.2000 75.1000 ;
	    RECT 2.2000 74.4000 2.6000 74.8000 ;
	    RECT 1.5000 73.4000 2.6000 73.7000 ;
	    RECT 2.2000 71.1000 2.6000 73.4000 ;
	    RECT 5.2000 72.5000 5.5000 75.8000 ;
	    RECT 10.3000 75.8000 10.6000 77.9000 ;
	    RECT 11.8000 77.1000 12.2000 79.9000 ;
	    RECT 13.4000 77.9000 13.8000 79.9000 ;
	    RECT 11.8000 76.8000 12.9000 77.1000 ;
	    RECT 11.8000 75.9000 12.2000 76.8000 ;
	    RECT 10.3000 75.5000 11.5000 75.8000 ;
	    RECT 5.8000 75.1000 6.6000 75.2000 ;
	    RECT 5.8000 74.8000 8.9000 75.1000 ;
	    RECT 10.2000 74.8000 10.6000 75.2000 ;
	    RECT 6.6000 73.8000 7.4000 74.2000 ;
	    RECT 8.6000 74.1000 8.9000 74.8000 ;
	    RECT 9.4000 74.1000 9.8000 74.6000 ;
	    RECT 10.3000 74.4000 10.6000 74.8000 ;
	    RECT 8.6000 73.8000 9.8000 74.1000 ;
	    RECT 10.2000 74.0000 10.8000 74.4000 ;
	    RECT 11.2000 73.8000 11.5000 75.5000 ;
	    RECT 11.9000 75.2000 12.2000 75.9000 ;
	    RECT 12.6000 76.2000 12.9000 76.8000 ;
	    RECT 12.6000 75.8000 13.0000 76.2000 ;
	    RECT 13.5000 75.8000 13.8000 77.9000 ;
	    RECT 15.0000 76.1000 15.4000 79.9000 ;
	    RECT 15.8000 76.8000 16.2000 77.2000 ;
	    RECT 15.8000 76.1000 16.1000 76.8000 ;
	    RECT 15.0000 75.8000 16.1000 76.1000 ;
	    RECT 13.5000 75.5000 14.7000 75.8000 ;
	    RECT 11.8000 74.8000 12.2000 75.2000 ;
	    RECT 13.4000 74.8000 13.8000 75.2000 ;
	    RECT 11.2000 73.7000 11.6000 73.8000 ;
	    RECT 10.1000 73.5000 11.6000 73.7000 ;
	    RECT 9.5000 73.4000 11.6000 73.5000 ;
	    RECT 9.5000 73.2000 10.4000 73.4000 ;
	    RECT 6.2000 73.1000 6.6000 73.2000 ;
	    RECT 7.3000 73.1000 8.2000 73.2000 ;
	    RECT 9.5000 73.1000 9.8000 73.2000 ;
	    RECT 11.9000 73.1000 12.2000 74.8000 ;
	    RECT 12.6000 73.8000 13.0000 74.6000 ;
	    RECT 13.5000 74.4000 13.8000 74.8000 ;
	    RECT 13.5000 74.1000 14.0000 74.4000 ;
	    RECT 13.6000 74.0000 14.0000 74.1000 ;
	    RECT 14.4000 73.8000 14.7000 75.5000 ;
	    RECT 15.1000 75.2000 15.4000 75.8000 ;
	    RECT 15.0000 74.8000 15.4000 75.2000 ;
	    RECT 14.4000 73.7000 14.8000 73.8000 ;
	    RECT 13.3000 73.5000 14.8000 73.7000 ;
	    RECT 12.7000 73.4000 14.8000 73.5000 ;
	    RECT 12.7000 73.2000 13.6000 73.4000 ;
	    RECT 12.7000 73.1000 13.0000 73.2000 ;
	    RECT 15.1000 73.1000 15.4000 74.8000 ;
	    RECT 15.8000 73.4000 16.2000 74.2000 ;
	    RECT 6.2000 72.8000 8.2000 73.1000 ;
	    RECT 5.2000 72.2000 7.2000 72.5000 ;
	    RECT 5.2000 72.1000 5.8000 72.2000 ;
	    RECT 5.4000 71.1000 5.8000 72.1000 ;
	    RECT 6.9000 71.8000 7.4000 72.2000 ;
	    RECT 7.0000 71.1000 7.4000 71.8000 ;
	    RECT 9.4000 71.1000 9.8000 73.1000 ;
	    RECT 11.5000 72.6000 12.2000 73.1000 ;
	    RECT 11.5000 71.1000 11.9000 72.6000 ;
	    RECT 12.6000 71.1000 13.0000 73.1000 ;
	    RECT 14.7000 72.6000 15.4000 73.1000 ;
	    RECT 16.6000 73.1000 17.0000 79.9000 ;
	    RECT 18.2000 77.9000 18.6000 79.9000 ;
	    RECT 18.3000 77.8000 18.6000 77.9000 ;
	    RECT 19.8000 77.9000 20.2000 79.9000 ;
	    RECT 19.8000 77.8000 20.1000 77.9000 ;
	    RECT 18.3000 77.5000 20.1000 77.8000 ;
	    RECT 17.4000 75.8000 17.8000 76.6000 ;
	    RECT 18.3000 76.2000 18.6000 77.5000 ;
	    RECT 19.0000 77.1000 19.4000 77.2000 ;
	    RECT 21.7000 77.1000 22.1000 79.9000 ;
	    RECT 19.0000 76.8000 22.1000 77.1000 ;
	    RECT 19.0000 76.4000 19.4000 76.8000 ;
	    RECT 21.7000 76.2000 22.1000 76.8000 ;
	    RECT 18.2000 75.8000 18.6000 76.2000 ;
	    RECT 18.3000 74.2000 18.6000 75.8000 ;
	    RECT 20.6000 75.4000 21.0000 76.2000 ;
	    RECT 21.4000 75.9000 22.1000 76.2000 ;
	    RECT 21.4000 75.2000 21.7000 75.9000 ;
	    RECT 23.8000 75.6000 24.2000 79.9000 ;
	    RECT 22.2000 75.4000 24.2000 75.6000 ;
	    RECT 22.1000 75.3000 24.2000 75.4000 ;
	    RECT 19.0000 74.8000 20.2000 75.2000 ;
	    RECT 21.4000 74.8000 21.8000 75.2000 ;
	    RECT 22.1000 75.0000 22.5000 75.3000 ;
	    RECT 18.3000 74.1000 19.1000 74.2000 ;
	    RECT 18.3000 73.9000 19.2000 74.1000 ;
	    RECT 16.6000 72.8000 17.5000 73.1000 ;
	    RECT 14.7000 71.1000 15.1000 72.6000 ;
	    RECT 17.1000 72.2000 17.5000 72.8000 ;
	    RECT 17.1000 71.8000 17.8000 72.2000 ;
	    RECT 17.1000 71.1000 17.5000 71.8000 ;
	    RECT 18.8000 71.1000 19.2000 73.9000 ;
	    RECT 21.4000 73.1000 21.7000 74.8000 ;
	    RECT 22.1000 73.5000 22.4000 75.0000 ;
	    RECT 22.8000 74.2000 23.2000 74.6000 ;
	    RECT 22.9000 73.8000 23.4000 74.2000 ;
	    RECT 22.1000 73.2000 23.3000 73.5000 ;
	    RECT 24.6000 73.4000 25.0000 74.2000 ;
	    RECT 21.4000 71.1000 21.8000 73.1000 ;
	    RECT 23.0000 72.1000 23.3000 73.2000 ;
	    RECT 23.8000 72.4000 24.2000 73.2000 ;
	    RECT 25.4000 73.1000 25.8000 79.9000 ;
	    RECT 26.2000 75.8000 26.6000 76.6000 ;
	    RECT 27.8000 76.4000 28.2000 79.9000 ;
	    RECT 27.7000 75.9000 28.2000 76.4000 ;
	    RECT 29.4000 76.2000 29.8000 79.9000 ;
	    RECT 31.5000 76.3000 31.9000 79.9000 ;
	    RECT 33.9000 79.2000 34.3000 79.9000 ;
	    RECT 33.9000 78.8000 34.6000 79.2000 ;
	    RECT 33.9000 76.3000 34.3000 78.8000 ;
	    RECT 28.5000 75.9000 29.8000 76.2000 ;
	    RECT 31.0000 75.9000 31.9000 76.3000 ;
	    RECT 33.4000 75.9000 34.3000 76.3000 ;
	    RECT 35.3000 76.2000 35.7000 79.9000 ;
	    RECT 35.0000 75.9000 35.7000 76.2000 ;
	    RECT 27.7000 74.2000 28.0000 75.9000 ;
	    RECT 28.5000 74.9000 28.8000 75.9000 ;
	    RECT 31.1000 75.2000 31.4000 75.9000 ;
	    RECT 28.3000 74.5000 28.8000 74.9000 ;
	    RECT 27.7000 73.8000 28.2000 74.2000 ;
	    RECT 27.7000 73.2000 28.0000 73.8000 ;
	    RECT 28.5000 73.7000 28.8000 74.5000 ;
	    RECT 29.3000 74.8000 29.8000 75.2000 ;
	    RECT 31.0000 74.8000 31.4000 75.2000 ;
	    RECT 31.8000 75.1000 32.2000 75.6000 ;
	    RECT 33.5000 75.1000 33.8000 75.9000 ;
	    RECT 31.8000 74.8000 33.8000 75.1000 ;
	    RECT 34.2000 75.1000 34.6000 75.6000 ;
	    RECT 35.0000 75.2000 35.3000 75.9000 ;
	    RECT 37.4000 75.6000 37.8000 79.9000 ;
	    RECT 38.5000 76.3000 38.9000 79.9000 ;
	    RECT 38.5000 75.9000 39.4000 76.3000 ;
	    RECT 39.0000 75.8000 39.4000 75.9000 ;
	    RECT 40.6000 75.8000 41.0000 76.6000 ;
	    RECT 35.8000 75.4000 37.8000 75.6000 ;
	    RECT 35.7000 75.3000 37.8000 75.4000 ;
	    RECT 35.0000 75.1000 35.4000 75.2000 ;
	    RECT 34.2000 74.8000 35.4000 75.1000 ;
	    RECT 35.7000 75.0000 36.1000 75.3000 ;
	    RECT 29.3000 74.4000 29.7000 74.8000 ;
	    RECT 31.1000 74.2000 31.4000 74.8000 ;
	    RECT 33.5000 74.2000 33.8000 74.8000 ;
	    RECT 31.0000 73.8000 31.4000 74.2000 ;
	    RECT 33.4000 73.8000 33.8000 74.2000 ;
	    RECT 28.5000 73.4000 29.8000 73.7000 ;
	    RECT 25.4000 72.8000 26.3000 73.1000 ;
	    RECT 27.7000 72.8000 28.2000 73.2000 ;
	    RECT 25.9000 72.2000 26.3000 72.8000 ;
	    RECT 23.0000 71.1000 23.4000 72.1000 ;
	    RECT 25.9000 71.8000 26.6000 72.2000 ;
	    RECT 25.9000 71.1000 26.3000 71.8000 ;
	    RECT 27.8000 71.1000 28.2000 72.8000 ;
	    RECT 29.4000 71.1000 29.8000 73.4000 ;
	    RECT 30.2000 72.4000 30.6000 73.2000 ;
	    RECT 31.1000 72.1000 31.4000 73.8000 ;
	    RECT 32.6000 72.4000 33.0000 73.2000 ;
	    RECT 33.5000 72.1000 33.8000 73.8000 ;
	    RECT 31.0000 71.1000 31.4000 72.1000 ;
	    RECT 33.4000 71.1000 33.8000 72.1000 ;
	    RECT 35.0000 73.1000 35.3000 74.8000 ;
	    RECT 35.7000 73.5000 36.0000 75.0000 ;
	    RECT 38.2000 74.8000 38.6000 75.6000 ;
	    RECT 36.4000 74.2000 36.8000 74.6000 ;
	    RECT 39.0000 74.2000 39.3000 75.8000 ;
	    RECT 36.5000 73.8000 37.0000 74.2000 ;
	    RECT 39.0000 73.8000 39.4000 74.2000 ;
	    RECT 40.6000 74.1000 41.0000 74.2000 ;
	    RECT 41.4000 74.1000 41.8000 79.9000 ;
	    RECT 43.3000 79.2000 43.7000 79.9000 ;
	    RECT 43.3000 78.8000 44.2000 79.2000 ;
	    RECT 43.3000 76.3000 43.7000 78.8000 ;
	    RECT 43.3000 75.9000 44.2000 76.3000 ;
	    RECT 43.0000 74.8000 43.4000 75.6000 ;
	    RECT 43.8000 74.2000 44.1000 75.9000 ;
	    RECT 40.6000 73.8000 41.8000 74.1000 ;
	    RECT 35.7000 73.2000 36.9000 73.5000 ;
	    RECT 35.0000 71.1000 35.4000 73.1000 ;
	    RECT 36.6000 72.1000 36.9000 73.2000 ;
	    RECT 37.4000 72.4000 37.8000 73.2000 ;
	    RECT 39.0000 72.1000 39.3000 73.8000 ;
	    RECT 39.8000 72.4000 40.2000 73.2000 ;
	    RECT 41.4000 73.1000 41.8000 73.8000 ;
	    RECT 42.2000 74.1000 42.6000 74.2000 ;
	    RECT 43.0000 74.1000 43.4000 74.2000 ;
	    RECT 42.2000 73.8000 43.4000 74.1000 ;
	    RECT 43.8000 73.8000 44.2000 74.2000 ;
	    RECT 42.2000 73.4000 42.6000 73.8000 ;
	    RECT 40.9000 72.8000 41.8000 73.1000 ;
	    RECT 36.6000 71.1000 37.0000 72.1000 ;
	    RECT 39.0000 71.1000 39.4000 72.1000 ;
	    RECT 40.9000 71.1000 41.3000 72.8000 ;
	    RECT 43.8000 72.1000 44.1000 73.8000 ;
	    RECT 45.4000 73.4000 45.8000 74.2000 ;
	    RECT 44.6000 72.4000 45.0000 73.2000 ;
	    RECT 46.2000 73.1000 46.6000 79.9000 ;
	    RECT 47.0000 76.1000 47.4000 76.6000 ;
	    RECT 49.4000 76.1000 49.8000 76.2000 ;
	    RECT 47.0000 75.8000 49.8000 76.1000 ;
	    RECT 50.2000 74.1000 50.6000 79.9000 ;
	    RECT 51.0000 76.2000 51.4000 79.9000 ;
	    RECT 52.6000 76.2000 53.0000 79.9000 ;
	    RECT 51.0000 75.9000 53.0000 76.2000 ;
	    RECT 53.4000 75.9000 53.8000 79.9000 ;
	    RECT 54.2000 75.9000 54.6000 79.9000 ;
	    RECT 55.0000 76.2000 55.4000 79.9000 ;
	    RECT 56.6000 76.2000 57.0000 79.9000 ;
	    RECT 55.0000 75.9000 57.0000 76.2000 ;
	    RECT 51.4000 75.2000 51.8000 75.4000 ;
	    RECT 53.4000 75.2000 53.7000 75.9000 ;
	    RECT 54.3000 75.2000 54.6000 75.9000 ;
	    RECT 58.2000 75.6000 58.6000 79.9000 ;
	    RECT 59.8000 75.6000 60.2000 79.9000 ;
	    RECT 56.2000 75.2000 56.6000 75.4000 ;
	    RECT 58.2000 75.2000 60.2000 75.6000 ;
	    RECT 51.0000 74.9000 51.8000 75.2000 ;
	    RECT 52.6000 74.9000 53.8000 75.2000 ;
	    RECT 51.0000 74.8000 51.4000 74.9000 ;
	    RECT 51.0000 74.1000 51.4000 74.2000 ;
	    RECT 50.2000 73.8000 51.4000 74.1000 ;
	    RECT 51.8000 73.8000 52.2000 74.6000 ;
	    RECT 46.2000 72.8000 47.1000 73.1000 ;
	    RECT 46.7000 72.1000 47.1000 72.8000 ;
	    RECT 49.4000 72.4000 49.8000 73.2000 ;
	    RECT 47.8000 72.1000 48.2000 72.2000 ;
	    RECT 43.8000 71.1000 44.2000 72.1000 ;
	    RECT 46.7000 71.8000 48.2000 72.1000 ;
	    RECT 46.7000 71.1000 47.1000 71.8000 ;
	    RECT 50.2000 71.1000 50.6000 73.8000 ;
	    RECT 52.6000 73.1000 52.9000 74.9000 ;
	    RECT 53.4000 74.8000 53.8000 74.9000 ;
	    RECT 54.2000 74.9000 55.4000 75.2000 ;
	    RECT 56.2000 75.1000 57.0000 75.2000 ;
	    RECT 58.2000 75.1000 58.6000 75.2000 ;
	    RECT 56.2000 74.9000 58.6000 75.1000 ;
	    RECT 54.2000 74.8000 54.6000 74.9000 ;
	    RECT 53.4000 73.1000 53.8000 73.2000 ;
	    RECT 54.2000 73.1000 54.6000 73.2000 ;
	    RECT 55.1000 73.1000 55.4000 74.9000 ;
	    RECT 56.6000 74.8000 58.6000 74.9000 ;
	    RECT 55.8000 73.8000 56.2000 74.6000 ;
	    RECT 56.6000 74.2000 56.9000 74.8000 ;
	    RECT 56.6000 73.8000 57.0000 74.2000 ;
	    RECT 57.4000 73.4000 57.8000 74.2000 ;
	    RECT 59.8000 73.8000 60.2000 75.2000 ;
	    RECT 58.2000 73.4000 60.2000 73.8000 ;
	    RECT 52.6000 71.1000 53.0000 73.1000 ;
	    RECT 53.4000 72.8000 54.6000 73.1000 ;
	    RECT 53.3000 72.4000 53.7000 72.8000 ;
	    RECT 54.3000 72.4000 54.7000 72.8000 ;
	    RECT 55.0000 71.1000 55.4000 73.1000 ;
	    RECT 58.2000 71.1000 58.6000 73.4000 ;
	    RECT 59.8000 71.1000 60.2000 73.4000 ;
	    RECT 61.4000 75.6000 61.8000 79.9000 ;
	    RECT 63.5000 77.9000 64.1000 79.9000 ;
	    RECT 65.8000 77.9000 66.2000 79.9000 ;
	    RECT 68.0000 78.2000 68.4000 79.9000 ;
	    RECT 68.0000 77.9000 69.0000 78.2000 ;
	    RECT 63.8000 77.5000 64.2000 77.9000 ;
	    RECT 65.9000 77.6000 66.2000 77.9000 ;
	    RECT 65.5000 77.3000 67.3000 77.6000 ;
	    RECT 68.6000 77.5000 69.0000 77.9000 ;
	    RECT 65.5000 77.2000 65.9000 77.3000 ;
	    RECT 66.9000 77.2000 67.3000 77.3000 ;
	    RECT 63.4000 76.6000 64.1000 77.0000 ;
	    RECT 63.8000 76.1000 64.1000 76.6000 ;
	    RECT 64.9000 76.5000 66.0000 76.8000 ;
	    RECT 64.9000 76.4000 65.3000 76.5000 ;
	    RECT 63.8000 75.8000 65.0000 76.1000 ;
	    RECT 61.4000 75.3000 63.5000 75.6000 ;
	    RECT 61.4000 73.6000 61.8000 75.3000 ;
	    RECT 63.1000 75.2000 63.5000 75.3000 ;
	    RECT 62.3000 74.9000 62.7000 75.0000 ;
	    RECT 62.3000 74.6000 64.2000 74.9000 ;
	    RECT 63.8000 74.5000 64.2000 74.6000 ;
	    RECT 64.7000 74.2000 65.0000 75.8000 ;
	    RECT 65.7000 75.9000 66.0000 76.5000 ;
	    RECT 66.3000 76.5000 66.7000 76.6000 ;
	    RECT 68.6000 76.5000 69.0000 76.6000 ;
	    RECT 66.3000 76.2000 69.0000 76.5000 ;
	    RECT 65.7000 75.7000 68.1000 75.9000 ;
	    RECT 70.2000 75.7000 70.6000 79.9000 ;
	    RECT 71.0000 76.2000 71.4000 79.9000 ;
	    RECT 73.2000 79.2000 74.0000 79.9000 ;
	    RECT 73.2000 78.8000 74.6000 79.2000 ;
	    RECT 71.8000 76.2000 72.2000 76.3000 ;
	    RECT 73.2000 76.2000 74.0000 78.8000 ;
	    RECT 71.0000 75.9000 72.2000 76.2000 ;
	    RECT 73.0000 75.9000 74.0000 76.2000 ;
	    RECT 75.1000 76.2000 75.5000 76.3000 ;
	    RECT 75.8000 76.2000 76.2000 79.9000 ;
	    RECT 75.1000 75.9000 76.2000 76.2000 ;
	    RECT 76.9000 76.3000 77.3000 79.9000 ;
	    RECT 76.9000 75.9000 77.8000 76.3000 ;
	    RECT 65.7000 75.6000 70.6000 75.7000 ;
	    RECT 67.7000 75.5000 70.6000 75.6000 ;
	    RECT 67.8000 75.4000 70.6000 75.5000 ;
	    RECT 73.0000 75.2000 73.3000 75.9000 ;
	    RECT 75.1000 75.6000 75.4000 75.9000 ;
	    RECT 73.7000 75.3000 75.4000 75.6000 ;
	    RECT 73.7000 75.2000 74.1000 75.3000 ;
	    RECT 67.0000 75.1000 67.4000 75.2000 ;
	    RECT 67.0000 74.8000 69.5000 75.1000 ;
	    RECT 72.6000 74.9000 73.3000 75.2000 ;
	    RECT 74.8000 74.9000 75.2000 75.0000 ;
	    RECT 72.6000 74.8000 73.5000 74.9000 ;
	    RECT 67.8000 74.7000 68.2000 74.8000 ;
	    RECT 69.1000 74.7000 69.5000 74.8000 ;
	    RECT 73.0000 74.6000 73.5000 74.8000 ;
	    RECT 68.3000 74.2000 68.7000 74.3000 ;
	    RECT 64.7000 73.9000 70.2000 74.2000 ;
	    RECT 64.9000 73.8000 65.3000 73.9000 ;
	    RECT 61.4000 73.3000 63.3000 73.6000 ;
	    RECT 61.4000 71.1000 61.8000 73.3000 ;
	    RECT 62.9000 73.2000 63.3000 73.3000 ;
	    RECT 67.8000 72.8000 68.1000 73.9000 ;
	    RECT 69.4000 73.8000 70.2000 73.9000 ;
	    RECT 71.0000 73.8000 71.8000 74.2000 ;
	    RECT 72.4000 73.8000 72.8000 74.2000 ;
	    RECT 72.5000 73.6000 72.8000 73.8000 ;
	    RECT 66.9000 72.7000 67.3000 72.8000 ;
	    RECT 63.8000 72.1000 64.2000 72.5000 ;
	    RECT 65.9000 72.4000 67.3000 72.7000 ;
	    RECT 67.8000 72.4000 68.2000 72.8000 ;
	    RECT 65.9000 72.1000 66.2000 72.4000 ;
	    RECT 68.6000 72.1000 69.0000 72.5000 ;
	    RECT 63.5000 71.8000 64.2000 72.1000 ;
	    RECT 63.5000 71.1000 64.1000 71.8000 ;
	    RECT 65.8000 71.1000 66.2000 72.1000 ;
	    RECT 68.0000 71.8000 69.0000 72.1000 ;
	    RECT 68.0000 71.1000 68.4000 71.8000 ;
	    RECT 70.2000 71.1000 70.6000 73.5000 ;
	    RECT 71.8000 73.4000 72.2000 73.5000 ;
	    RECT 71.0000 73.1000 72.2000 73.4000 ;
	    RECT 72.5000 73.2000 72.9000 73.6000 ;
	    RECT 71.0000 71.1000 71.4000 73.1000 ;
	    RECT 73.2000 72.9000 73.5000 74.6000 ;
	    RECT 73.9000 74.6000 75.2000 74.9000 ;
	    RECT 76.6000 74.8000 77.0000 75.6000 ;
	    RECT 73.9000 74.3000 74.2000 74.6000 ;
	    RECT 73.8000 73.9000 74.2000 74.3000 ;
	    RECT 77.4000 74.2000 77.7000 75.9000 ;
	    RECT 75.4000 74.1000 76.2000 74.2000 ;
	    RECT 77.4000 74.1000 77.8000 74.2000 ;
	    RECT 74.5000 73.8000 77.8000 74.1000 ;
	    RECT 74.5000 73.6000 74.8000 73.8000 ;
	    RECT 73.8000 73.3000 74.8000 73.6000 ;
	    RECT 75.1000 73.4000 75.5000 73.5000 ;
	    RECT 73.8000 73.2000 74.6000 73.3000 ;
	    RECT 75.1000 73.1000 76.2000 73.4000 ;
	    RECT 73.2000 71.1000 74.0000 72.9000 ;
	    RECT 75.8000 71.1000 76.2000 73.1000 ;
	    RECT 77.4000 72.1000 77.7000 73.8000 ;
	    RECT 79.0000 73.4000 79.4000 74.2000 ;
	    RECT 78.2000 72.4000 78.6000 73.2000 ;
	    RECT 79.8000 73.1000 80.2000 79.9000 ;
	    RECT 80.6000 75.8000 81.0000 76.6000 ;
	    RECT 81.4000 75.8000 81.8000 79.9000 ;
	    RECT 83.0000 77.9000 83.4000 79.9000 ;
	    RECT 85.4000 77.9000 85.8000 79.9000 ;
	    RECT 83.0000 75.8000 83.3000 77.9000 ;
	    RECT 85.5000 77.8000 85.8000 77.9000 ;
	    RECT 87.0000 77.9000 87.4000 79.9000 ;
	    RECT 87.8000 77.9000 88.2000 79.9000 ;
	    RECT 87.0000 77.8000 87.3000 77.9000 ;
	    RECT 85.5000 77.5000 87.3000 77.8000 ;
	    RECT 86.2000 76.4000 86.6000 77.2000 ;
	    RECT 87.0000 76.2000 87.3000 77.5000 ;
	    RECT 87.9000 77.8000 88.2000 77.9000 ;
	    RECT 89.4000 77.8000 89.8000 79.9000 ;
	    RECT 87.9000 77.5000 89.7000 77.8000 ;
	    RECT 91.0000 77.5000 91.4000 79.5000 ;
	    RECT 93.1000 79.2000 93.5000 79.9000 ;
	    RECT 93.1000 78.8000 93.8000 79.2000 ;
	    RECT 87.9000 76.2000 88.2000 77.5000 ;
	    RECT 88.6000 76.4000 89.0000 77.2000 ;
	    RECT 81.4000 75.2000 81.7000 75.8000 ;
	    RECT 82.1000 75.5000 83.3000 75.8000 ;
	    RECT 81.4000 74.8000 81.8000 75.2000 ;
	    RECT 81.4000 73.1000 81.7000 74.8000 ;
	    RECT 82.1000 73.8000 82.4000 75.5000 ;
	    RECT 84.6000 75.4000 85.0000 76.2000 ;
	    RECT 87.0000 75.8000 87.4000 76.2000 ;
	    RECT 87.8000 75.8000 88.2000 76.2000 ;
	    RECT 83.0000 74.8000 83.4000 75.2000 ;
	    RECT 85.4000 74.8000 86.2000 75.2000 ;
	    RECT 83.0000 74.4000 83.3000 74.8000 ;
	    RECT 82.8000 74.1000 83.3000 74.4000 ;
	    RECT 82.8000 74.0000 83.2000 74.1000 ;
	    RECT 83.8000 73.8000 84.2000 74.6000 ;
	    RECT 87.0000 74.2000 87.3000 75.8000 ;
	    RECT 86.5000 74.1000 87.3000 74.2000 ;
	    RECT 86.4000 73.9000 87.3000 74.1000 ;
	    RECT 87.9000 74.2000 88.2000 75.8000 ;
	    RECT 90.2000 75.4000 90.6000 76.2000 ;
	    RECT 91.0000 75.8000 91.3000 77.5000 ;
	    RECT 93.1000 76.4000 93.5000 78.8000 ;
	    RECT 96.6000 77.9000 97.0000 79.9000 ;
	    RECT 96.7000 77.8000 97.0000 77.9000 ;
	    RECT 98.2000 77.9000 98.6000 79.9000 ;
	    RECT 100.7000 79.6000 102.5000 79.9000 ;
	    RECT 100.7000 79.5000 101.0000 79.6000 ;
	    RECT 98.2000 77.8000 98.5000 77.9000 ;
	    RECT 96.7000 77.5000 98.5000 77.8000 ;
	    RECT 97.4000 76.4000 97.8000 77.2000 ;
	    RECT 93.1000 76.1000 93.9000 76.4000 ;
	    RECT 98.2000 76.2000 98.5000 77.5000 ;
	    RECT 100.6000 76.5000 101.0000 79.5000 ;
	    RECT 102.2000 79.5000 102.5000 79.6000 ;
	    RECT 103.0000 79.6000 105.0000 79.9000 ;
	    RECT 101.4000 76.5000 101.8000 79.3000 ;
	    RECT 102.2000 76.7000 102.6000 79.5000 ;
	    RECT 103.0000 77.0000 103.4000 79.6000 ;
	    RECT 103.8000 76.9000 104.2000 79.3000 ;
	    RECT 104.6000 76.9000 105.0000 79.6000 ;
	    RECT 103.8000 76.7000 104.1000 76.9000 ;
	    RECT 102.2000 76.5000 104.1000 76.7000 ;
	    RECT 101.5000 76.2000 101.8000 76.5000 ;
	    RECT 102.3000 76.4000 104.1000 76.5000 ;
	    RECT 104.7000 76.6000 105.0000 76.9000 ;
	    RECT 106.2000 76.9000 106.6000 79.9000 ;
	    RECT 107.0000 77.9000 107.4000 79.9000 ;
	    RECT 107.1000 77.8000 107.4000 77.9000 ;
	    RECT 108.6000 77.9000 109.0000 79.9000 ;
	    RECT 108.6000 77.8000 108.9000 77.9000 ;
	    RECT 107.1000 77.5000 108.9000 77.8000 ;
	    RECT 106.2000 76.6000 106.5000 76.9000 ;
	    RECT 104.7000 76.3000 106.5000 76.6000 ;
	    RECT 107.1000 76.2000 107.4000 77.5000 ;
	    RECT 108.6000 77.2000 108.9000 77.5000 ;
	    RECT 107.8000 76.4000 108.2000 77.2000 ;
	    RECT 108.6000 76.8000 109.0000 77.2000 ;
	    RECT 111.5000 76.2000 111.9000 79.9000 ;
	    RECT 114.7000 77.2000 115.1000 79.9000 ;
	    RECT 112.2000 76.8000 112.6000 77.2000 ;
	    RECT 114.2000 76.8000 115.1000 77.2000 ;
	    RECT 115.4000 76.8000 115.8000 77.2000 ;
	    RECT 112.3000 76.2000 112.6000 76.8000 ;
	    RECT 114.7000 76.2000 115.1000 76.8000 ;
	    RECT 115.5000 76.2000 115.8000 76.8000 ;
	    RECT 91.0000 75.5000 92.9000 75.8000 ;
	    RECT 89.0000 74.8000 89.8000 75.2000 ;
	    RECT 91.0000 74.4000 91.4000 75.2000 ;
	    RECT 91.8000 74.4000 92.2000 75.2000 ;
	    RECT 92.6000 74.5000 92.9000 75.5000 ;
	    RECT 87.9000 74.1000 88.7000 74.2000 ;
	    RECT 92.6000 74.1000 93.3000 74.5000 ;
	    RECT 93.6000 74.2000 93.9000 76.1000 ;
	    RECT 94.2000 74.8000 94.6000 75.6000 ;
	    RECT 95.8000 75.4000 96.2000 76.2000 ;
	    RECT 98.2000 75.8000 98.6000 76.2000 ;
	    RECT 99.0000 76.1000 99.4000 76.2000 ;
	    RECT 101.4000 76.1000 101.8000 76.2000 ;
	    RECT 99.0000 75.8000 103.1000 76.1000 ;
	    RECT 107.0000 75.8000 107.4000 76.2000 ;
	    RECT 96.6000 74.8000 97.4000 75.2000 ;
	    RECT 98.2000 74.2000 98.5000 75.8000 ;
	    RECT 87.9000 73.9000 88.8000 74.1000 ;
	    RECT 92.6000 73.9000 93.1000 74.1000 ;
	    RECT 82.0000 73.7000 82.4000 73.8000 ;
	    RECT 82.0000 73.5000 83.5000 73.7000 ;
	    RECT 82.0000 73.4000 84.1000 73.5000 ;
	    RECT 83.2000 73.2000 84.1000 73.4000 ;
	    RECT 83.8000 73.1000 84.1000 73.2000 ;
	    RECT 79.8000 72.8000 80.7000 73.1000 ;
	    RECT 80.3000 72.2000 80.7000 72.8000 ;
	    RECT 81.4000 72.6000 82.1000 73.1000 ;
	    RECT 77.4000 71.1000 77.8000 72.1000 ;
	    RECT 79.8000 71.8000 80.7000 72.2000 ;
	    RECT 80.3000 71.1000 80.7000 71.8000 ;
	    RECT 81.7000 71.1000 82.1000 72.6000 ;
	    RECT 83.8000 71.1000 84.2000 73.1000 ;
	    RECT 86.4000 71.1000 86.8000 73.9000 ;
	    RECT 88.4000 71.1000 88.8000 73.9000 ;
	    RECT 91.0000 73.6000 93.1000 73.9000 ;
	    RECT 93.6000 73.8000 94.6000 74.2000 ;
	    RECT 97.7000 74.1000 98.5000 74.2000 ;
	    RECT 97.6000 73.9000 98.5000 74.1000 ;
	    RECT 91.0000 72.5000 91.3000 73.6000 ;
	    RECT 93.6000 73.5000 93.9000 73.8000 ;
	    RECT 93.5000 73.3000 93.9000 73.5000 ;
	    RECT 93.1000 73.0000 93.9000 73.3000 ;
	    RECT 91.0000 71.5000 91.4000 72.5000 ;
	    RECT 93.1000 71.5000 93.5000 73.0000 ;
	    RECT 97.6000 71.1000 98.0000 73.9000 ;
	    RECT 102.8000 72.5000 103.1000 75.8000 ;
	    RECT 103.4000 74.8000 104.2000 75.2000 ;
	    RECT 107.1000 74.2000 107.4000 75.8000 ;
	    RECT 108.2000 74.8000 109.0000 75.2000 ;
	    RECT 109.4000 75.1000 109.8000 76.2000 ;
	    RECT 111.5000 75.9000 112.0000 76.2000 ;
	    RECT 112.3000 75.9000 113.0000 76.2000 ;
	    RECT 114.7000 75.9000 115.2000 76.2000 ;
	    RECT 115.5000 75.9000 116.2000 76.2000 ;
	    RECT 116.6000 75.9000 117.0000 79.9000 ;
	    RECT 117.4000 76.2000 117.8000 79.9000 ;
	    RECT 119.0000 76.2000 119.4000 79.9000 ;
	    RECT 120.6000 77.9000 121.0000 79.9000 ;
	    RECT 117.4000 75.9000 119.4000 76.2000 ;
	    RECT 111.7000 75.2000 112.0000 75.9000 ;
	    RECT 112.6000 75.8000 113.0000 75.9000 ;
	    RECT 111.0000 75.1000 111.4000 75.2000 ;
	    RECT 109.4000 74.8000 111.4000 75.1000 ;
	    RECT 111.0000 74.4000 111.4000 74.8000 ;
	    RECT 111.7000 74.8000 112.2000 75.2000 ;
	    RECT 111.7000 74.2000 112.0000 74.8000 ;
	    RECT 114.2000 74.4000 114.6000 75.2000 ;
	    RECT 114.9000 74.2000 115.2000 75.9000 ;
	    RECT 115.8000 75.8000 116.2000 75.9000 ;
	    RECT 116.7000 75.2000 117.0000 75.9000 ;
	    RECT 120.7000 75.8000 121.0000 77.9000 ;
	    RECT 122.2000 75.9000 122.6000 79.9000 ;
	    RECT 124.3000 76.2000 124.7000 79.9000 ;
	    RECT 127.0000 77.9000 127.4000 79.9000 ;
	    RECT 125.0000 76.8000 125.4000 77.2000 ;
	    RECT 125.1000 76.2000 125.4000 76.8000 ;
	    RECT 124.3000 75.9000 124.8000 76.2000 ;
	    RECT 125.1000 75.9000 125.8000 76.2000 ;
	    RECT 120.7000 75.5000 121.9000 75.8000 ;
	    RECT 118.6000 75.2000 119.0000 75.4000 ;
	    RECT 116.6000 74.9000 117.8000 75.2000 ;
	    RECT 118.6000 74.9000 119.4000 75.2000 ;
	    RECT 116.6000 74.8000 117.0000 74.9000 ;
	    RECT 104.2000 74.1000 105.0000 74.2000 ;
	    RECT 106.2000 74.1000 106.6000 74.2000 ;
	    RECT 104.2000 73.8000 106.6000 74.1000 ;
	    RECT 107.1000 74.1000 107.9000 74.2000 ;
	    RECT 110.2000 74.1000 110.6000 74.2000 ;
	    RECT 107.1000 73.9000 108.0000 74.1000 ;
	    RECT 104.9000 72.8000 105.8000 73.2000 ;
	    RECT 102.8000 72.2000 104.8000 72.5000 ;
	    RECT 102.8000 72.1000 103.4000 72.2000 ;
	    RECT 103.0000 71.1000 103.4000 72.1000 ;
	    RECT 104.5000 72.1000 104.8000 72.2000 ;
	    RECT 104.5000 71.8000 105.0000 72.1000 ;
	    RECT 104.6000 71.1000 105.0000 71.8000 ;
	    RECT 107.6000 71.1000 108.0000 73.9000 ;
	    RECT 110.2000 73.8000 111.0000 74.1000 ;
	    RECT 111.7000 73.8000 113.0000 74.2000 ;
	    RECT 113.4000 74.1000 113.8000 74.2000 ;
	    RECT 113.4000 73.8000 114.2000 74.1000 ;
	    RECT 114.9000 73.8000 116.2000 74.2000 ;
	    RECT 110.6000 73.6000 111.0000 73.8000 ;
	    RECT 110.3000 73.1000 112.1000 73.3000 ;
	    RECT 112.6000 73.1000 112.9000 73.8000 ;
	    RECT 113.8000 73.6000 114.2000 73.8000 ;
	    RECT 113.5000 73.1000 115.3000 73.3000 ;
	    RECT 115.8000 73.1000 116.1000 73.8000 ;
	    RECT 110.2000 73.0000 112.2000 73.1000 ;
	    RECT 110.2000 71.1000 110.6000 73.0000 ;
	    RECT 111.8000 71.1000 112.2000 73.0000 ;
	    RECT 112.6000 71.1000 113.0000 73.1000 ;
	    RECT 113.4000 73.0000 115.4000 73.1000 ;
	    RECT 113.4000 71.1000 113.8000 73.0000 ;
	    RECT 115.0000 71.1000 115.4000 73.0000 ;
	    RECT 115.8000 71.1000 116.2000 73.1000 ;
	    RECT 116.6000 72.8000 117.0000 73.2000 ;
	    RECT 117.5000 73.1000 117.8000 74.9000 ;
	    RECT 119.0000 74.8000 119.4000 74.9000 ;
	    RECT 120.6000 74.8000 121.0000 75.2000 ;
	    RECT 118.2000 73.8000 118.6000 74.6000 ;
	    RECT 119.8000 73.8000 120.2000 74.6000 ;
	    RECT 120.7000 74.4000 121.0000 74.8000 ;
	    RECT 120.7000 74.1000 121.2000 74.4000 ;
	    RECT 120.8000 74.0000 121.2000 74.1000 ;
	    RECT 121.6000 73.8000 121.9000 75.5000 ;
	    RECT 122.3000 75.2000 122.6000 75.9000 ;
	    RECT 124.4000 75.8000 124.8000 75.9000 ;
	    RECT 125.4000 75.8000 125.8000 75.9000 ;
	    RECT 127.1000 75.8000 127.4000 77.9000 ;
	    RECT 128.6000 75.9000 129.0000 79.9000 ;
	    RECT 130.7000 79.2000 131.1000 79.9000 ;
	    RECT 130.2000 78.8000 131.1000 79.2000 ;
	    RECT 130.7000 76.2000 131.1000 78.8000 ;
	    RECT 131.4000 76.8000 131.8000 77.2000 ;
	    RECT 131.5000 76.2000 131.8000 76.8000 ;
	    RECT 130.7000 75.9000 131.2000 76.2000 ;
	    RECT 131.5000 75.9000 132.2000 76.2000 ;
	    RECT 122.2000 74.8000 122.6000 75.2000 ;
	    RECT 123.0000 75.1000 123.4000 75.2000 ;
	    RECT 123.8000 75.1000 124.2000 75.2000 ;
	    RECT 123.0000 74.8000 124.2000 75.1000 ;
	    RECT 121.6000 73.7000 122.0000 73.8000 ;
	    RECT 120.5000 73.5000 122.0000 73.7000 ;
	    RECT 119.9000 73.4000 122.0000 73.5000 ;
	    RECT 119.9000 73.2000 120.8000 73.4000 ;
	    RECT 119.9000 73.1000 120.2000 73.2000 ;
	    RECT 122.3000 73.1000 122.6000 74.8000 ;
	    RECT 123.8000 74.4000 124.2000 74.8000 ;
	    RECT 124.5000 74.2000 124.8000 75.8000 ;
	    RECT 127.1000 75.5000 128.3000 75.8000 ;
	    RECT 127.0000 74.8000 127.4000 75.2000 ;
	    RECT 123.0000 74.1000 123.4000 74.2000 ;
	    RECT 123.0000 73.8000 123.8000 74.1000 ;
	    RECT 124.5000 73.8000 125.8000 74.2000 ;
	    RECT 126.2000 73.8000 126.6000 74.6000 ;
	    RECT 127.1000 74.4000 127.4000 74.8000 ;
	    RECT 127.1000 74.1000 127.6000 74.4000 ;
	    RECT 127.2000 74.0000 127.6000 74.1000 ;
	    RECT 128.0000 73.8000 128.3000 75.5000 ;
	    RECT 128.7000 75.2000 129.0000 75.9000 ;
	    RECT 128.6000 75.1000 129.0000 75.2000 ;
	    RECT 128.6000 74.8000 129.7000 75.1000 ;
	    RECT 123.4000 73.6000 123.8000 73.8000 ;
	    RECT 123.1000 73.1000 124.9000 73.3000 ;
	    RECT 125.4000 73.1000 125.7000 73.8000 ;
	    RECT 128.0000 73.7000 128.4000 73.8000 ;
	    RECT 126.9000 73.5000 128.4000 73.7000 ;
	    RECT 126.3000 73.4000 128.4000 73.5000 ;
	    RECT 126.3000 73.2000 127.2000 73.4000 ;
	    RECT 126.3000 73.1000 126.6000 73.2000 ;
	    RECT 128.7000 73.1000 129.0000 74.8000 ;
	    RECT 129.4000 74.2000 129.7000 74.8000 ;
	    RECT 130.2000 74.4000 130.6000 75.2000 ;
	    RECT 130.9000 74.2000 131.2000 75.9000 ;
	    RECT 131.8000 75.8000 132.2000 75.9000 ;
	    RECT 129.4000 74.1000 129.8000 74.2000 ;
	    RECT 129.4000 73.8000 130.2000 74.1000 ;
	    RECT 130.9000 73.8000 132.2000 74.2000 ;
	    RECT 129.8000 73.6000 130.2000 73.8000 ;
	    RECT 129.5000 73.1000 131.3000 73.3000 ;
	    RECT 131.8000 73.1000 132.1000 73.8000 ;
	    RECT 132.6000 73.4000 133.0000 74.2000 ;
	    RECT 116.7000 72.4000 117.1000 72.8000 ;
	    RECT 117.4000 71.1000 117.8000 73.1000 ;
	    RECT 119.8000 71.1000 120.2000 73.1000 ;
	    RECT 121.9000 72.6000 122.6000 73.1000 ;
	    RECT 123.0000 73.0000 125.0000 73.1000 ;
	    RECT 121.9000 72.2000 122.3000 72.6000 ;
	    RECT 121.9000 71.8000 122.6000 72.2000 ;
	    RECT 121.9000 71.1000 122.3000 71.8000 ;
	    RECT 123.0000 71.1000 123.4000 73.0000 ;
	    RECT 124.6000 71.1000 125.0000 73.0000 ;
	    RECT 125.4000 71.1000 125.8000 73.1000 ;
	    RECT 126.2000 71.1000 126.6000 73.1000 ;
	    RECT 128.3000 72.6000 129.0000 73.1000 ;
	    RECT 129.4000 73.0000 131.4000 73.1000 ;
	    RECT 128.3000 71.1000 128.7000 72.6000 ;
	    RECT 129.4000 71.1000 129.8000 73.0000 ;
	    RECT 131.0000 71.1000 131.4000 73.0000 ;
	    RECT 131.8000 71.1000 132.2000 73.1000 ;
	    RECT 133.4000 71.1000 133.8000 79.9000 ;
	    RECT 135.5000 76.2000 135.9000 79.9000 ;
	    RECT 138.7000 77.2000 139.1000 79.9000 ;
	    RECT 136.2000 76.8000 136.6000 77.2000 ;
	    RECT 138.2000 76.8000 139.1000 77.2000 ;
	    RECT 139.4000 76.8000 139.8000 77.2000 ;
	    RECT 136.3000 76.2000 136.6000 76.8000 ;
	    RECT 138.7000 76.2000 139.1000 76.8000 ;
	    RECT 139.5000 76.2000 139.8000 76.8000 ;
	    RECT 135.5000 75.9000 136.0000 76.2000 ;
	    RECT 136.3000 75.9000 137.0000 76.2000 ;
	    RECT 138.7000 75.9000 139.2000 76.2000 ;
	    RECT 139.5000 76.1000 140.2000 76.2000 ;
	    RECT 140.6000 76.1000 141.0000 79.9000 ;
	    RECT 139.5000 75.9000 141.0000 76.1000 ;
	    RECT 141.4000 76.2000 141.8000 79.9000 ;
	    RECT 143.0000 76.2000 143.4000 79.9000 ;
	    RECT 141.4000 75.9000 143.4000 76.2000 ;
	    RECT 143.8000 76.2000 144.2000 79.9000 ;
	    RECT 143.8000 75.9000 144.9000 76.2000 ;
	    RECT 135.0000 74.4000 135.4000 75.2000 ;
	    RECT 135.7000 74.2000 136.0000 75.9000 ;
	    RECT 136.6000 75.8000 137.0000 75.9000 ;
	    RECT 138.2000 74.4000 138.6000 75.2000 ;
	    RECT 138.9000 74.2000 139.2000 75.9000 ;
	    RECT 139.8000 75.8000 141.0000 75.9000 ;
	    RECT 140.7000 75.2000 141.0000 75.8000 ;
	    RECT 144.6000 75.6000 144.9000 75.9000 ;
	    RECT 142.6000 75.2000 143.0000 75.4000 ;
	    RECT 144.6000 75.2000 145.2000 75.6000 ;
	    RECT 140.6000 74.9000 141.8000 75.2000 ;
	    RECT 142.6000 74.9000 143.4000 75.2000 ;
	    RECT 140.6000 74.8000 141.0000 74.9000 ;
	    RECT 134.2000 74.1000 134.6000 74.2000 ;
	    RECT 135.7000 74.1000 137.0000 74.2000 ;
	    RECT 137.4000 74.1000 137.8000 74.2000 ;
	    RECT 134.2000 73.8000 135.0000 74.1000 ;
	    RECT 135.7000 73.8000 138.2000 74.1000 ;
	    RECT 138.9000 73.8000 140.2000 74.2000 ;
	    RECT 134.6000 73.6000 135.0000 73.8000 ;
	    RECT 134.3000 73.1000 136.1000 73.3000 ;
	    RECT 136.6000 73.1000 136.9000 73.8000 ;
	    RECT 137.8000 73.6000 138.2000 73.8000 ;
	    RECT 137.5000 73.1000 139.3000 73.3000 ;
	    RECT 139.8000 73.1000 140.1000 73.8000 ;
	    RECT 134.2000 73.0000 136.2000 73.1000 ;
	    RECT 134.2000 71.1000 134.6000 73.0000 ;
	    RECT 135.8000 71.1000 136.2000 73.0000 ;
	    RECT 136.6000 71.1000 137.0000 73.1000 ;
	    RECT 137.4000 73.0000 139.4000 73.1000 ;
	    RECT 137.4000 71.1000 137.8000 73.0000 ;
	    RECT 139.0000 71.1000 139.4000 73.0000 ;
	    RECT 139.8000 71.1000 140.2000 73.1000 ;
	    RECT 140.6000 72.8000 141.0000 73.2000 ;
	    RECT 141.5000 73.1000 141.8000 74.9000 ;
	    RECT 143.0000 74.8000 143.4000 74.9000 ;
	    RECT 142.2000 73.8000 142.6000 74.6000 ;
	    RECT 143.8000 74.4000 144.2000 75.2000 ;
	    RECT 144.6000 73.7000 144.9000 75.2000 ;
	    RECT 140.7000 72.4000 141.1000 72.8000 ;
	    RECT 141.4000 71.1000 141.8000 73.1000 ;
	    RECT 143.8000 73.4000 144.9000 73.7000 ;
	    RECT 143.8000 71.1000 144.2000 73.4000 ;
	    RECT 2.2000 67.6000 2.6000 69.9000 ;
	    RECT 1.5000 67.3000 2.6000 67.6000 ;
	    RECT 3.0000 67.7000 3.4000 69.9000 ;
	    RECT 5.1000 69.2000 5.7000 69.9000 ;
	    RECT 5.1000 68.9000 5.8000 69.2000 ;
	    RECT 7.4000 68.9000 7.8000 69.9000 ;
	    RECT 9.6000 69.2000 10.0000 69.9000 ;
	    RECT 9.6000 68.9000 10.6000 69.2000 ;
	    RECT 5.4000 68.5000 5.8000 68.9000 ;
	    RECT 7.5000 68.6000 7.8000 68.9000 ;
	    RECT 7.5000 68.3000 8.9000 68.6000 ;
	    RECT 8.5000 68.2000 8.9000 68.3000 ;
	    RECT 9.4000 68.2000 9.8000 68.6000 ;
	    RECT 10.2000 68.5000 10.6000 68.9000 ;
	    RECT 4.5000 67.7000 4.9000 67.8000 ;
	    RECT 3.0000 67.4000 5.0000 67.7000 ;
	    RECT 1.5000 65.8000 1.8000 67.3000 ;
	    RECT 2.2000 66.1000 2.6000 66.6000 ;
	    RECT 3.0000 66.1000 3.4000 67.4000 ;
	    RECT 4.6000 66.8000 5.0000 67.4000 ;
	    RECT 6.5000 67.1000 6.9000 67.2000 ;
	    RECT 9.4000 67.1000 9.7000 68.2000 ;
	    RECT 11.8000 67.5000 12.2000 69.9000 ;
	    RECT 11.0000 67.1000 11.8000 67.2000 ;
	    RECT 6.3000 66.8000 11.8000 67.1000 ;
	    RECT 12.6000 66.8000 13.0000 67.6000 ;
	    RECT 13.4000 67.1000 13.8000 69.9000 ;
	    RECT 14.2000 67.9000 14.6000 69.9000 ;
	    RECT 16.4000 68.1000 17.2000 69.9000 ;
	    RECT 14.2000 67.6000 15.4000 67.9000 ;
	    RECT 15.0000 67.5000 15.4000 67.6000 ;
	    RECT 15.7000 67.4000 16.1000 67.8000 ;
	    RECT 15.7000 67.2000 16.0000 67.4000 ;
	    RECT 14.2000 67.1000 15.0000 67.2000 ;
	    RECT 13.4000 66.8000 15.0000 67.1000 ;
	    RECT 15.6000 66.8000 16.0000 67.2000 ;
	    RECT 5.4000 66.4000 5.8000 66.5000 ;
	    RECT 2.2000 65.8000 3.4000 66.1000 ;
	    RECT 3.9000 66.1000 5.8000 66.4000 ;
	    RECT 3.9000 66.0000 4.3000 66.1000 ;
	    RECT 1.2000 65.4000 1.8000 65.8000 ;
	    RECT 1.5000 65.1000 1.8000 65.4000 ;
	    RECT 3.0000 65.7000 3.4000 65.8000 ;
	    RECT 4.7000 65.7000 5.1000 65.8000 ;
	    RECT 3.0000 65.4000 5.1000 65.7000 ;
	    RECT 1.5000 64.8000 2.6000 65.1000 ;
	    RECT 2.2000 61.1000 2.6000 64.8000 ;
	    RECT 3.0000 61.1000 3.4000 65.4000 ;
	    RECT 6.3000 65.2000 6.6000 66.8000 ;
	    RECT 9.9000 66.7000 10.3000 66.8000 ;
	    RECT 9.4000 66.2000 9.8000 66.3000 ;
	    RECT 10.7000 66.2000 11.1000 66.3000 ;
	    RECT 8.6000 65.9000 11.1000 66.2000 ;
	    RECT 8.6000 65.8000 9.0000 65.9000 ;
	    RECT 9.4000 65.5000 12.2000 65.6000 ;
	    RECT 9.3000 65.4000 12.2000 65.5000 ;
	    RECT 5.4000 64.9000 6.6000 65.2000 ;
	    RECT 7.3000 65.3000 12.2000 65.4000 ;
	    RECT 7.3000 65.1000 9.7000 65.3000 ;
	    RECT 5.4000 64.4000 5.7000 64.9000 ;
	    RECT 5.0000 64.0000 5.7000 64.4000 ;
	    RECT 6.5000 64.5000 6.9000 64.6000 ;
	    RECT 7.3000 64.5000 7.6000 65.1000 ;
	    RECT 6.5000 64.2000 7.6000 64.5000 ;
	    RECT 7.9000 64.5000 10.6000 64.8000 ;
	    RECT 7.9000 64.4000 8.3000 64.5000 ;
	    RECT 10.2000 64.4000 10.6000 64.5000 ;
	    RECT 7.1000 63.7000 7.5000 63.8000 ;
	    RECT 8.5000 63.7000 8.9000 63.8000 ;
	    RECT 5.4000 63.1000 5.8000 63.5000 ;
	    RECT 7.1000 63.4000 8.9000 63.7000 ;
	    RECT 7.5000 63.1000 7.8000 63.4000 ;
	    RECT 10.2000 63.1000 10.6000 63.5000 ;
	    RECT 5.1000 61.1000 5.7000 63.1000 ;
	    RECT 7.4000 61.1000 7.8000 63.1000 ;
	    RECT 9.6000 62.8000 10.6000 63.1000 ;
	    RECT 9.6000 61.1000 10.0000 62.8000 ;
	    RECT 11.8000 61.1000 12.2000 65.3000 ;
	    RECT 13.4000 61.1000 13.8000 66.8000 ;
	    RECT 14.2000 66.2000 14.5000 66.8000 ;
	    RECT 16.4000 66.4000 16.7000 68.1000 ;
	    RECT 19.0000 67.9000 19.4000 69.9000 ;
	    RECT 17.0000 67.7000 17.8000 67.8000 ;
	    RECT 17.0000 67.4000 18.0000 67.7000 ;
	    RECT 18.3000 67.6000 19.4000 67.9000 ;
	    RECT 21.4000 67.8000 21.8000 69.9000 ;
	    RECT 22.1000 68.2000 22.5000 68.6000 ;
	    RECT 22.2000 68.1000 22.6000 68.2000 ;
	    RECT 23.0000 68.1000 23.4000 69.9000 ;
	    RECT 22.2000 67.8000 23.4000 68.1000 ;
	    RECT 23.8000 68.0000 24.2000 69.9000 ;
	    RECT 25.4000 68.0000 25.8000 69.9000 ;
	    RECT 23.8000 67.9000 25.8000 68.0000 ;
	    RECT 18.3000 67.5000 18.7000 67.6000 ;
	    RECT 17.7000 67.2000 18.0000 67.4000 ;
	    RECT 17.0000 66.7000 17.4000 67.1000 ;
	    RECT 17.7000 66.9000 19.4000 67.2000 ;
	    RECT 18.6000 66.8000 19.4000 66.9000 ;
	    RECT 16.2000 66.2000 16.7000 66.4000 ;
	    RECT 14.2000 65.8000 14.6000 66.2000 ;
	    RECT 15.8000 66.1000 16.7000 66.2000 ;
	    RECT 17.1000 66.4000 17.4000 66.7000 ;
	    RECT 20.6000 66.4000 21.0000 67.2000 ;
	    RECT 17.1000 66.1000 18.4000 66.4000 ;
	    RECT 15.8000 65.8000 16.5000 66.1000 ;
	    RECT 18.0000 66.0000 18.4000 66.1000 ;
	    RECT 19.8000 66.1000 20.2000 66.2000 ;
	    RECT 21.4000 66.1000 21.7000 67.8000 ;
	    RECT 23.1000 67.2000 23.4000 67.8000 ;
	    RECT 23.9000 67.7000 25.7000 67.9000 ;
	    RECT 25.0000 67.2000 25.4000 67.4000 ;
	    RECT 23.0000 66.8000 24.3000 67.2000 ;
	    RECT 25.0000 66.9000 25.8000 67.2000 ;
	    RECT 26.8000 67.1000 27.2000 69.9000 ;
	    RECT 29.4000 67.9000 29.8000 69.9000 ;
	    RECT 30.2000 68.0000 30.6000 69.9000 ;
	    RECT 31.8000 68.0000 32.2000 69.9000 ;
	    RECT 30.2000 67.9000 32.2000 68.0000 ;
	    RECT 29.5000 67.2000 29.8000 67.9000 ;
	    RECT 30.3000 67.7000 32.1000 67.9000 ;
	    RECT 31.4000 67.2000 31.8000 67.4000 ;
	    RECT 25.4000 66.8000 25.8000 66.9000 ;
	    RECT 26.3000 66.9000 27.2000 67.1000 ;
	    RECT 26.3000 66.8000 27.1000 66.9000 ;
	    RECT 29.4000 66.8000 30.7000 67.2000 ;
	    RECT 31.4000 66.9000 32.2000 67.2000 ;
	    RECT 34.4000 67.1000 34.8000 69.9000 ;
	    RECT 35.8000 67.9000 36.2000 69.9000 ;
	    RECT 36.6000 68.0000 37.0000 69.9000 ;
	    RECT 38.2000 68.0000 38.6000 69.9000 ;
	    RECT 36.6000 67.9000 38.6000 68.0000 ;
	    RECT 35.9000 67.2000 36.2000 67.9000 ;
	    RECT 36.7000 67.7000 38.5000 67.9000 ;
	    RECT 37.8000 67.2000 38.2000 67.4000 ;
	    RECT 34.4000 66.9000 35.3000 67.1000 ;
	    RECT 31.8000 66.8000 32.2000 66.9000 ;
	    RECT 34.5000 66.8000 35.3000 66.9000 ;
	    RECT 35.8000 66.8000 37.1000 67.2000 ;
	    RECT 37.8000 66.9000 38.6000 67.2000 ;
	    RECT 38.2000 66.8000 38.6000 66.9000 ;
	    RECT 22.2000 66.1000 22.6000 66.2000 ;
	    RECT 19.8000 65.8000 20.6000 66.1000 ;
	    RECT 21.4000 65.8000 22.6000 66.1000 ;
	    RECT 16.2000 65.1000 16.5000 65.8000 ;
	    RECT 16.9000 65.7000 17.3000 65.8000 ;
	    RECT 16.9000 65.4000 18.6000 65.7000 ;
	    RECT 20.2000 65.6000 20.6000 65.8000 ;
	    RECT 18.3000 65.1000 18.6000 65.4000 ;
	    RECT 22.2000 65.1000 22.5000 65.8000 ;
	    RECT 23.0000 65.1000 23.4000 65.2000 ;
	    RECT 24.0000 65.1000 24.3000 66.8000 ;
	    RECT 24.6000 65.8000 25.0000 66.6000 ;
	    RECT 26.3000 65.2000 26.6000 66.8000 ;
	    RECT 27.4000 65.8000 28.2000 66.2000 ;
	    RECT 14.2000 64.8000 15.4000 65.1000 ;
	    RECT 16.2000 64.8000 17.2000 65.1000 ;
	    RECT 14.2000 61.1000 14.6000 64.8000 ;
	    RECT 15.0000 64.7000 15.4000 64.8000 ;
	    RECT 16.4000 61.1000 17.2000 64.8000 ;
	    RECT 18.3000 64.8000 19.4000 65.1000 ;
	    RECT 18.3000 64.7000 18.7000 64.8000 ;
	    RECT 19.0000 61.1000 19.4000 64.8000 ;
	    RECT 19.8000 64.8000 21.8000 65.1000 ;
	    RECT 19.8000 61.1000 20.2000 64.8000 ;
	    RECT 21.4000 61.1000 21.8000 64.8000 ;
	    RECT 22.2000 61.1000 22.6000 65.1000 ;
	    RECT 23.0000 64.8000 23.7000 65.1000 ;
	    RECT 24.0000 64.8000 24.5000 65.1000 ;
	    RECT 26.2000 64.8000 26.6000 65.2000 ;
	    RECT 28.6000 64.8000 29.0000 65.6000 ;
	    RECT 29.4000 65.1000 29.8000 65.2000 ;
	    RECT 30.4000 65.1000 30.7000 66.8000 ;
	    RECT 31.0000 65.8000 31.4000 66.6000 ;
	    RECT 33.4000 65.8000 34.2000 66.2000 ;
	    RECT 29.4000 64.8000 30.1000 65.1000 ;
	    RECT 30.4000 64.8000 30.9000 65.1000 ;
	    RECT 32.6000 64.8000 33.0000 65.6000 ;
	    RECT 35.0000 65.2000 35.3000 66.8000 ;
	    RECT 36.8000 65.2000 37.1000 66.8000 ;
	    RECT 37.4000 66.1000 37.8000 66.6000 ;
	    RECT 39.0000 66.1000 39.4000 69.9000 ;
	    RECT 40.9000 69.2000 41.3000 69.9000 ;
	    RECT 40.6000 68.8000 41.3000 69.2000 ;
	    RECT 39.8000 67.8000 40.2000 68.6000 ;
	    RECT 40.9000 68.2000 41.3000 68.8000 ;
	    RECT 44.3000 68.2000 44.7000 69.9000 ;
	    RECT 45.5000 68.2000 45.9000 68.6000 ;
	    RECT 40.9000 67.9000 41.8000 68.2000 ;
	    RECT 37.4000 65.8000 39.4000 66.1000 ;
	    RECT 35.0000 64.8000 35.4000 65.2000 ;
	    RECT 35.8000 65.1000 36.2000 65.2000 ;
	    RECT 35.8000 64.8000 36.5000 65.1000 ;
	    RECT 36.8000 64.8000 37.8000 65.2000 ;
	    RECT 23.4000 64.2000 23.7000 64.8000 ;
	    RECT 23.4000 63.8000 23.8000 64.2000 ;
	    RECT 24.1000 61.1000 24.5000 64.8000 ;
	    RECT 26.3000 63.5000 26.6000 64.8000 ;
	    RECT 27.0000 63.8000 27.4000 64.6000 ;
	    RECT 29.8000 64.2000 30.1000 64.8000 ;
	    RECT 29.8000 64.1000 30.2000 64.2000 ;
	    RECT 27.8000 63.8000 30.2000 64.1000 ;
	    RECT 27.8000 63.5000 28.1000 63.8000 ;
	    RECT 26.3000 63.2000 28.1000 63.5000 ;
	    RECT 26.3000 63.1000 26.6000 63.2000 ;
	    RECT 26.2000 61.1000 26.6000 63.1000 ;
	    RECT 27.8000 63.1000 28.1000 63.2000 ;
	    RECT 27.8000 61.1000 28.2000 63.1000 ;
	    RECT 30.5000 62.2000 30.9000 64.8000 ;
	    RECT 34.2000 63.8000 34.6000 64.6000 ;
	    RECT 35.0000 64.2000 35.3000 64.8000 ;
	    RECT 36.2000 64.2000 36.5000 64.8000 ;
	    RECT 35.0000 63.8000 35.4000 64.2000 ;
	    RECT 36.2000 63.8000 36.6000 64.2000 ;
	    RECT 35.0000 63.5000 35.3000 63.8000 ;
	    RECT 33.5000 63.2000 35.3000 63.5000 ;
	    RECT 33.5000 63.1000 33.8000 63.2000 ;
	    RECT 30.5000 61.8000 31.4000 62.2000 ;
	    RECT 30.5000 61.1000 30.9000 61.8000 ;
	    RECT 33.4000 61.1000 33.8000 63.1000 ;
	    RECT 35.0000 63.1000 35.3000 63.2000 ;
	    RECT 35.0000 61.1000 35.4000 63.1000 ;
	    RECT 36.9000 61.1000 37.3000 64.8000 ;
	    RECT 39.0000 61.1000 39.4000 65.8000 ;
	    RECT 40.6000 64.4000 41.0000 65.2000 ;
	    RECT 41.4000 61.1000 41.8000 67.9000 ;
	    RECT 43.8000 67.9000 44.7000 68.2000 ;
	    RECT 42.2000 66.8000 42.6000 67.6000 ;
	    RECT 43.0000 66.8000 43.4000 67.6000 ;
	    RECT 43.8000 61.1000 44.2000 67.9000 ;
	    RECT 45.4000 67.8000 45.8000 68.2000 ;
	    RECT 46.2000 67.9000 46.6000 69.9000 ;
	    RECT 52.6000 68.9000 53.0000 69.9000 ;
	    RECT 54.2000 69.2000 54.6000 69.9000 ;
	    RECT 45.4000 66.1000 45.8000 66.2000 ;
	    RECT 46.3000 66.1000 46.6000 67.9000 ;
	    RECT 52.4000 68.8000 53.0000 68.9000 ;
	    RECT 54.1000 68.8000 54.6000 69.2000 ;
	    RECT 52.4000 68.5000 54.4000 68.8000 ;
	    RECT 47.0000 66.4000 47.4000 67.2000 ;
	    RECT 47.8000 66.1000 48.2000 66.2000 ;
	    RECT 48.6000 66.1000 49.0000 66.2000 ;
	    RECT 45.4000 65.8000 46.6000 66.1000 ;
	    RECT 47.4000 65.8000 49.0000 66.1000 ;
	    RECT 44.6000 65.1000 45.0000 65.2000 ;
	    RECT 45.5000 65.1000 45.8000 65.8000 ;
	    RECT 47.4000 65.6000 47.8000 65.8000 ;
	    RECT 52.4000 65.2000 52.7000 68.5000 ;
	    RECT 54.5000 67.8000 55.4000 68.2000 ;
	    RECT 56.6000 68.0000 57.0000 69.9000 ;
	    RECT 58.2000 68.0000 58.6000 69.9000 ;
	    RECT 56.6000 67.9000 58.6000 68.0000 ;
	    RECT 59.0000 67.9000 59.4000 69.9000 ;
	    RECT 61.1000 68.2000 61.5000 69.9000 ;
	    RECT 63.0000 68.2000 63.4000 69.9000 ;
	    RECT 60.6000 67.9000 61.5000 68.2000 ;
	    RECT 62.9000 67.9000 63.4000 68.2000 ;
	    RECT 56.7000 67.7000 58.5000 67.9000 ;
	    RECT 57.0000 67.2000 57.4000 67.4000 ;
	    RECT 59.0000 67.2000 59.3000 67.9000 ;
	    RECT 53.8000 66.8000 54.6000 67.2000 ;
	    RECT 55.8000 67.1000 56.2000 67.2000 ;
	    RECT 56.6000 67.1000 57.4000 67.2000 ;
	    RECT 55.8000 66.9000 57.4000 67.1000 ;
	    RECT 58.1000 67.1000 59.4000 67.2000 ;
	    RECT 59.8000 67.1000 60.2000 67.6000 ;
	    RECT 55.8000 66.8000 57.0000 66.9000 ;
	    RECT 58.1000 66.8000 60.2000 67.1000 ;
	    RECT 60.6000 67.1000 61.0000 67.9000 ;
	    RECT 62.9000 67.2000 63.2000 67.9000 ;
	    RECT 64.6000 67.6000 65.0000 69.9000 ;
	    RECT 65.4000 67.9000 65.8000 69.9000 ;
	    RECT 67.6000 68.1000 68.4000 69.9000 ;
	    RECT 65.4000 67.6000 66.5000 67.9000 ;
	    RECT 67.0000 67.7000 67.8000 67.8000 ;
	    RECT 63.7000 67.3000 65.0000 67.6000 ;
	    RECT 66.1000 67.5000 66.5000 67.6000 ;
	    RECT 66.8000 67.4000 67.8000 67.7000 ;
	    RECT 61.4000 67.1000 61.8000 67.2000 ;
	    RECT 60.6000 66.8000 61.8000 67.1000 ;
	    RECT 62.9000 66.8000 63.4000 67.2000 ;
	    RECT 53.0000 65.8000 53.8000 66.2000 ;
	    RECT 55.0000 66.1000 55.4000 66.2000 ;
	    RECT 56.6000 66.1000 57.0000 66.2000 ;
	    RECT 57.4000 66.1000 57.8000 66.6000 ;
	    RECT 55.0000 65.8000 57.8000 66.1000 ;
	    RECT 44.6000 64.8000 45.8000 65.1000 ;
	    RECT 44.6000 64.4000 45.0000 64.8000 ;
	    RECT 45.4000 61.1000 45.8000 64.8000 ;
	    RECT 46.2000 64.8000 48.2000 65.1000 ;
	    RECT 51.0000 64.9000 52.7000 65.2000 ;
	    RECT 58.1000 65.1000 58.4000 66.8000 ;
	    RECT 59.0000 65.1000 59.4000 65.2000 ;
	    RECT 51.0000 64.8000 51.4000 64.9000 ;
	    RECT 46.2000 61.1000 46.6000 64.8000 ;
	    RECT 47.8000 61.1000 48.2000 64.8000 ;
	    RECT 51.1000 64.5000 51.4000 64.8000 ;
	    RECT 57.9000 64.8000 58.4000 65.1000 ;
	    RECT 58.7000 64.8000 59.4000 65.1000 ;
	    RECT 51.9000 64.5000 53.7000 64.6000 ;
	    RECT 50.2000 61.5000 50.6000 64.5000 ;
	    RECT 51.0000 61.7000 51.4000 64.5000 ;
	    RECT 51.8000 64.3000 53.7000 64.5000 ;
	    RECT 50.3000 61.4000 50.6000 61.5000 ;
	    RECT 51.8000 61.5000 52.2000 64.3000 ;
	    RECT 53.4000 64.1000 53.7000 64.3000 ;
	    RECT 54.3000 64.4000 56.1000 64.7000 ;
	    RECT 54.3000 64.1000 54.6000 64.4000 ;
	    RECT 51.8000 61.4000 52.1000 61.5000 ;
	    RECT 50.3000 61.1000 52.1000 61.4000 ;
	    RECT 52.6000 61.4000 53.0000 64.0000 ;
	    RECT 53.4000 61.7000 53.8000 64.1000 ;
	    RECT 54.2000 61.4000 54.6000 64.1000 ;
	    RECT 52.6000 61.1000 54.6000 61.4000 ;
	    RECT 55.8000 64.1000 56.1000 64.4000 ;
	    RECT 55.8000 61.1000 56.2000 64.1000 ;
	    RECT 57.9000 61.1000 58.3000 64.8000 ;
	    RECT 58.7000 64.2000 59.0000 64.8000 ;
	    RECT 58.6000 63.8000 59.0000 64.2000 ;
	    RECT 60.6000 61.1000 61.0000 66.8000 ;
	    RECT 62.9000 65.2000 63.2000 66.8000 ;
	    RECT 63.7000 66.5000 64.0000 67.3000 ;
	    RECT 66.8000 67.2000 67.1000 67.4000 ;
	    RECT 65.4000 66.9000 67.1000 67.2000 ;
	    RECT 65.4000 66.8000 66.2000 66.9000 ;
	    RECT 67.4000 66.7000 67.8000 67.1000 ;
	    RECT 63.5000 66.1000 64.0000 66.5000 ;
	    RECT 61.4000 64.4000 61.8000 65.2000 ;
	    RECT 62.9000 64.6000 63.4000 65.2000 ;
	    RECT 63.7000 65.1000 64.0000 66.1000 ;
	    RECT 64.5000 66.2000 64.9000 66.6000 ;
	    RECT 67.4000 66.4000 67.7000 66.7000 ;
	    RECT 64.5000 65.8000 65.0000 66.2000 ;
	    RECT 66.4000 66.1000 67.7000 66.4000 ;
	    RECT 68.1000 66.4000 68.4000 68.1000 ;
	    RECT 70.2000 67.9000 70.6000 69.9000 ;
	    RECT 68.7000 67.4000 69.1000 67.8000 ;
	    RECT 69.4000 67.6000 70.6000 67.9000 ;
	    RECT 71.0000 67.6000 71.4000 69.9000 ;
	    RECT 72.6000 68.2000 73.0000 69.9000 ;
	    RECT 76.6000 68.9000 77.0000 69.9000 ;
	    RECT 78.2000 69.2000 78.6000 69.9000 ;
	    RECT 76.4000 68.8000 77.0000 68.9000 ;
	    RECT 78.1000 68.8000 78.6000 69.2000 ;
	    RECT 81.4000 68.8000 81.8000 69.9000 ;
	    RECT 83.3000 69.2000 83.7000 69.9000 ;
	    RECT 83.0000 68.8000 83.7000 69.2000 ;
	    RECT 76.4000 68.5000 78.4000 68.8000 ;
	    RECT 72.6000 67.9000 73.1000 68.2000 ;
	    RECT 69.4000 67.5000 69.8000 67.6000 ;
	    RECT 68.8000 67.2000 69.1000 67.4000 ;
	    RECT 71.0000 67.3000 72.3000 67.6000 ;
	    RECT 68.8000 66.8000 69.2000 67.2000 ;
	    RECT 69.8000 66.8000 70.6000 67.2000 ;
	    RECT 68.1000 66.2000 68.6000 66.4000 ;
	    RECT 71.1000 66.2000 71.5000 66.6000 ;
	    RECT 68.1000 66.1000 69.0000 66.2000 ;
	    RECT 66.4000 66.0000 66.8000 66.1000 ;
	    RECT 68.3000 65.8000 69.0000 66.1000 ;
	    RECT 70.2000 66.1000 70.6000 66.2000 ;
	    RECT 71.0000 66.1000 71.5000 66.2000 ;
	    RECT 70.2000 65.8000 71.5000 66.1000 ;
	    RECT 72.0000 66.5000 72.3000 67.3000 ;
	    RECT 72.8000 67.2000 73.1000 67.9000 ;
	    RECT 72.6000 66.8000 73.1000 67.2000 ;
	    RECT 72.0000 66.1000 72.5000 66.5000 ;
	    RECT 67.5000 65.7000 67.9000 65.8000 ;
	    RECT 66.2000 65.4000 67.9000 65.7000 ;
	    RECT 66.2000 65.1000 66.5000 65.4000 ;
	    RECT 68.3000 65.1000 68.6000 65.8000 ;
	    RECT 72.0000 65.1000 72.3000 66.1000 ;
	    RECT 72.8000 65.1000 73.1000 66.8000 ;
	    RECT 76.4000 65.2000 76.7000 68.5000 ;
	    RECT 78.5000 67.8000 79.4000 68.2000 ;
	    RECT 81.4000 67.2000 81.7000 68.8000 ;
	    RECT 82.2000 67.8000 82.6000 68.6000 ;
	    RECT 83.3000 68.4000 83.7000 68.8000 ;
	    RECT 83.0000 67.9000 83.7000 68.4000 ;
	    RECT 85.4000 67.9000 85.8000 69.9000 ;
	    RECT 87.5000 69.2000 87.9000 69.9000 ;
	    RECT 87.5000 68.8000 88.2000 69.2000 ;
	    RECT 87.5000 68.2000 87.9000 68.8000 ;
	    RECT 89.9000 68.2000 90.3000 69.9000 ;
	    RECT 91.8000 68.9000 92.2000 69.9000 ;
	    RECT 95.0000 69.2000 95.4000 69.9000 ;
	    RECT 95.0000 68.9000 95.5000 69.2000 ;
	    RECT 87.0000 67.9000 87.9000 68.2000 ;
	    RECT 89.4000 68.1000 90.3000 68.2000 ;
	    RECT 91.0000 68.1000 91.4000 68.6000 ;
	    RECT 77.8000 67.1000 78.6000 67.2000 ;
	    RECT 80.6000 67.1000 81.0000 67.2000 ;
	    RECT 77.8000 66.8000 81.0000 67.1000 ;
	    RECT 81.4000 66.8000 81.8000 67.2000 ;
	    RECT 77.0000 65.8000 77.8000 66.2000 ;
	    RECT 80.6000 65.4000 81.0000 66.2000 ;
	    RECT 63.7000 64.8000 65.0000 65.1000 ;
	    RECT 63.0000 61.1000 63.4000 64.6000 ;
	    RECT 64.6000 61.1000 65.0000 64.8000 ;
	    RECT 65.4000 64.8000 66.5000 65.1000 ;
	    RECT 65.4000 61.1000 65.8000 64.8000 ;
	    RECT 66.1000 64.7000 66.5000 64.8000 ;
	    RECT 67.6000 64.8000 68.6000 65.1000 ;
	    RECT 69.4000 64.8000 70.6000 65.1000 ;
	    RECT 67.6000 61.1000 68.4000 64.8000 ;
	    RECT 69.4000 64.7000 69.8000 64.8000 ;
	    RECT 70.2000 61.1000 70.6000 64.8000 ;
	    RECT 71.0000 64.8000 72.3000 65.1000 ;
	    RECT 71.0000 61.1000 71.4000 64.8000 ;
	    RECT 72.6000 64.6000 73.1000 65.1000 ;
	    RECT 75.0000 64.9000 76.7000 65.2000 ;
	    RECT 81.4000 65.1000 81.7000 66.8000 ;
	    RECT 83.0000 66.2000 83.3000 67.9000 ;
	    RECT 85.4000 67.8000 85.7000 67.9000 ;
	    RECT 84.8000 67.6000 85.7000 67.8000 ;
	    RECT 83.6000 67.5000 85.7000 67.6000 ;
	    RECT 83.6000 67.3000 85.1000 67.5000 ;
	    RECT 83.6000 67.2000 84.0000 67.3000 ;
	    RECT 83.0000 65.8000 83.4000 66.2000 ;
	    RECT 83.0000 65.1000 83.3000 65.8000 ;
	    RECT 83.7000 65.5000 84.0000 67.2000 ;
	    RECT 84.4000 66.9000 84.8000 67.0000 ;
	    RECT 84.4000 66.6000 84.9000 66.9000 ;
	    RECT 84.6000 66.2000 84.9000 66.6000 ;
	    RECT 85.4000 66.4000 85.8000 67.2000 ;
	    RECT 86.2000 66.8000 86.6000 67.6000 ;
	    RECT 84.6000 65.8000 85.0000 66.2000 ;
	    RECT 83.7000 65.2000 84.9000 65.5000 ;
	    RECT 75.0000 64.8000 75.4000 64.9000 ;
	    RECT 72.6000 61.1000 73.0000 64.6000 ;
	    RECT 75.1000 64.5000 75.4000 64.8000 ;
	    RECT 80.9000 64.7000 81.8000 65.1000 ;
	    RECT 75.9000 64.5000 77.7000 64.6000 ;
	    RECT 74.2000 61.5000 74.6000 64.5000 ;
	    RECT 75.0000 61.7000 75.4000 64.5000 ;
	    RECT 75.8000 64.3000 77.7000 64.5000 ;
	    RECT 74.3000 61.4000 74.6000 61.5000 ;
	    RECT 75.8000 61.5000 76.2000 64.3000 ;
	    RECT 77.4000 64.1000 77.7000 64.3000 ;
	    RECT 78.3000 64.4000 80.1000 64.7000 ;
	    RECT 78.3000 64.1000 78.6000 64.4000 ;
	    RECT 75.8000 61.4000 76.1000 61.5000 ;
	    RECT 74.3000 61.1000 76.1000 61.4000 ;
	    RECT 76.6000 61.4000 77.0000 64.0000 ;
	    RECT 77.4000 61.7000 77.8000 64.1000 ;
	    RECT 78.2000 61.4000 78.6000 64.1000 ;
	    RECT 76.6000 61.1000 78.6000 61.4000 ;
	    RECT 79.8000 64.1000 80.1000 64.4000 ;
	    RECT 79.8000 61.1000 80.2000 64.1000 ;
	    RECT 80.9000 61.1000 81.3000 64.7000 ;
	    RECT 83.0000 61.1000 83.4000 65.1000 ;
	    RECT 84.6000 63.1000 84.9000 65.2000 ;
	    RECT 84.6000 61.1000 85.0000 63.1000 ;
	    RECT 87.0000 61.1000 87.4000 67.9000 ;
	    RECT 89.4000 67.8000 91.4000 68.1000 ;
	    RECT 88.6000 66.8000 89.0000 67.6000 ;
	    RECT 87.8000 64.4000 88.2000 65.2000 ;
	    RECT 89.4000 61.1000 89.8000 67.8000 ;
	    RECT 91.9000 67.2000 92.2000 68.9000 ;
	    RECT 95.2000 68.8000 95.5000 68.9000 ;
	    RECT 96.6000 69.1000 97.0000 69.9000 ;
	    RECT 99.8000 69.1000 100.2000 69.2000 ;
	    RECT 101.7000 69.1000 102.1000 69.9000 ;
	    RECT 96.6000 68.8000 100.2000 69.1000 ;
	    RECT 100.6000 68.8000 102.1000 69.1000 ;
	    RECT 95.2000 68.5000 97.2000 68.8000 ;
	    RECT 94.2000 67.8000 95.1000 68.2000 ;
	    RECT 91.8000 66.8000 92.2000 67.2000 ;
	    RECT 92.6000 67.1000 93.0000 67.2000 ;
	    RECT 95.0000 67.1000 95.8000 67.2000 ;
	    RECT 92.6000 66.8000 95.8000 67.1000 ;
	    RECT 91.0000 66.1000 91.4000 66.2000 ;
	    RECT 91.9000 66.1000 92.2000 66.8000 ;
	    RECT 91.0000 65.8000 92.2000 66.1000 ;
	    RECT 90.2000 64.4000 90.6000 65.2000 ;
	    RECT 91.9000 65.1000 92.2000 65.8000 ;
	    RECT 92.6000 65.4000 93.0000 66.2000 ;
	    RECT 95.8000 65.8000 96.6000 66.2000 ;
	    RECT 96.9000 65.2000 97.2000 68.5000 ;
	    RECT 100.6000 68.2000 100.9000 68.8000 ;
	    RECT 101.7000 68.4000 102.1000 68.8000 ;
	    RECT 100.6000 67.8000 101.0000 68.2000 ;
	    RECT 101.4000 67.9000 102.1000 68.4000 ;
	    RECT 103.8000 67.9000 104.2000 69.9000 ;
	    RECT 104.9000 68.2000 105.3000 69.9000 ;
	    RECT 104.9000 67.9000 105.8000 68.2000 ;
	    RECT 101.4000 66.2000 101.7000 67.9000 ;
	    RECT 103.8000 67.8000 104.1000 67.9000 ;
	    RECT 103.2000 67.6000 104.1000 67.8000 ;
	    RECT 102.0000 67.5000 104.1000 67.6000 ;
	    RECT 102.0000 67.3000 103.5000 67.5000 ;
	    RECT 102.0000 67.2000 102.4000 67.3000 ;
	    RECT 101.4000 65.8000 101.8000 66.2000 ;
	    RECT 91.8000 64.7000 92.7000 65.1000 ;
	    RECT 96.9000 64.9000 98.6000 65.2000 ;
	    RECT 98.2000 64.8000 98.6000 64.9000 ;
	    RECT 101.4000 65.1000 101.7000 65.8000 ;
	    RECT 102.1000 65.5000 102.4000 67.2000 ;
	    RECT 103.8000 67.1000 104.2000 67.2000 ;
	    RECT 104.6000 67.1000 105.0000 67.2000 ;
	    RECT 102.8000 66.9000 103.2000 67.0000 ;
	    RECT 102.8000 66.6000 103.3000 66.9000 ;
	    RECT 103.0000 66.2000 103.3000 66.6000 ;
	    RECT 103.8000 66.8000 105.0000 67.1000 ;
	    RECT 103.8000 66.4000 104.2000 66.8000 ;
	    RECT 103.0000 65.8000 103.4000 66.2000 ;
	    RECT 104.6000 66.1000 105.0000 66.2000 ;
	    RECT 105.4000 66.1000 105.8000 67.9000 ;
	    RECT 106.2000 66.8000 106.6000 67.6000 ;
	    RECT 107.6000 67.1000 108.0000 69.9000 ;
	    RECT 110.2000 68.0000 110.6000 69.9000 ;
	    RECT 111.8000 68.0000 112.2000 69.9000 ;
	    RECT 110.2000 67.9000 112.2000 68.0000 ;
	    RECT 112.6000 67.9000 113.0000 69.9000 ;
	    RECT 114.0000 69.1000 114.4000 69.9000 ;
	    RECT 115.0000 69.1000 115.4000 69.2000 ;
	    RECT 114.0000 68.8000 115.4000 69.1000 ;
	    RECT 117.4000 68.9000 117.8000 69.9000 ;
	    RECT 110.3000 67.7000 112.1000 67.9000 ;
	    RECT 110.6000 67.2000 111.0000 67.4000 ;
	    RECT 112.6000 67.2000 112.9000 67.9000 ;
	    RECT 107.1000 66.9000 108.0000 67.1000 ;
	    RECT 110.2000 66.9000 111.0000 67.2000 ;
	    RECT 107.1000 66.8000 107.9000 66.9000 ;
	    RECT 110.2000 66.8000 110.6000 66.9000 ;
	    RECT 111.7000 66.8000 113.0000 67.2000 ;
	    RECT 114.0000 67.1000 114.4000 68.8000 ;
	    RECT 116.6000 67.8000 117.0000 68.6000 ;
	    RECT 117.5000 67.2000 117.8000 68.9000 ;
	    RECT 113.5000 66.9000 114.4000 67.1000 ;
	    RECT 113.5000 66.8000 114.3000 66.9000 ;
	    RECT 117.4000 66.8000 117.8000 67.2000 ;
	    RECT 120.8000 67.1000 121.2000 69.9000 ;
	    RECT 122.2000 68.0000 122.6000 69.9000 ;
	    RECT 123.8000 68.0000 124.2000 69.9000 ;
	    RECT 122.2000 67.9000 124.2000 68.0000 ;
	    RECT 122.3000 67.7000 124.1000 67.9000 ;
	    RECT 124.6000 67.8000 125.0000 69.9000 ;
	    RECT 122.6000 67.2000 123.0000 67.4000 ;
	    RECT 124.6000 67.2000 124.9000 67.8000 ;
	    RECT 120.8000 66.9000 121.7000 67.1000 ;
	    RECT 120.9000 66.8000 121.7000 66.9000 ;
	    RECT 122.2000 66.9000 123.0000 67.2000 ;
	    RECT 122.2000 66.8000 122.6000 66.9000 ;
	    RECT 123.7000 66.8000 125.0000 67.2000 ;
	    RECT 104.6000 65.8000 105.8000 66.1000 ;
	    RECT 102.1000 65.2000 103.3000 65.5000 ;
	    RECT 92.3000 61.1000 92.7000 64.7000 ;
	    RECT 93.5000 64.4000 95.3000 64.7000 ;
	    RECT 93.5000 64.1000 93.8000 64.4000 ;
	    RECT 93.4000 61.1000 93.8000 64.1000 ;
	    RECT 95.0000 64.1000 95.3000 64.4000 ;
	    RECT 95.9000 64.5000 97.7000 64.6000 ;
	    RECT 98.2000 64.5000 98.5000 64.8000 ;
	    RECT 95.9000 64.3000 97.8000 64.5000 ;
	    RECT 95.9000 64.1000 96.2000 64.3000 ;
	    RECT 95.0000 61.4000 95.4000 64.1000 ;
	    RECT 95.8000 61.7000 96.2000 64.1000 ;
	    RECT 96.6000 61.4000 97.0000 64.0000 ;
	    RECT 97.4000 61.5000 97.8000 64.3000 ;
	    RECT 98.2000 61.7000 98.6000 64.5000 ;
	    RECT 95.0000 61.1000 97.0000 61.4000 ;
	    RECT 97.5000 61.4000 97.8000 61.5000 ;
	    RECT 99.0000 61.5000 99.4000 64.5000 ;
	    RECT 99.0000 61.4000 99.3000 61.5000 ;
	    RECT 97.5000 61.1000 99.3000 61.4000 ;
	    RECT 101.4000 61.1000 101.8000 65.1000 ;
	    RECT 103.0000 63.1000 103.3000 65.2000 ;
	    RECT 103.8000 65.1000 104.2000 65.2000 ;
	    RECT 104.6000 65.1000 105.0000 65.2000 ;
	    RECT 103.8000 64.8000 105.0000 65.1000 ;
	    RECT 104.6000 64.4000 105.0000 64.8000 ;
	    RECT 103.0000 61.1000 103.4000 63.1000 ;
	    RECT 105.4000 61.1000 105.8000 65.8000 ;
	    RECT 107.1000 65.2000 107.4000 66.8000 ;
	    RECT 108.2000 65.8000 109.0000 66.2000 ;
	    RECT 111.0000 65.8000 111.4000 66.6000 ;
	    RECT 107.0000 64.8000 107.4000 65.2000 ;
	    RECT 109.4000 64.8000 109.8000 65.6000 ;
	    RECT 111.7000 65.1000 112.0000 66.8000 ;
	    RECT 113.5000 65.2000 113.8000 66.8000 ;
	    RECT 114.6000 65.8000 115.4000 66.2000 ;
	    RECT 112.6000 65.1000 113.0000 65.2000 ;
	    RECT 111.5000 64.8000 112.0000 65.1000 ;
	    RECT 112.3000 64.8000 113.0000 65.1000 ;
	    RECT 113.4000 64.8000 113.8000 65.2000 ;
	    RECT 115.8000 64.8000 116.2000 65.6000 ;
	    RECT 117.5000 65.2000 117.8000 66.8000 ;
	    RECT 118.2000 65.4000 118.6000 66.2000 ;
	    RECT 119.8000 65.8000 120.6000 66.2000 ;
	    RECT 117.4000 65.1000 117.8000 65.2000 ;
	    RECT 106.2000 64.1000 106.6000 64.2000 ;
	    RECT 107.1000 64.1000 107.4000 64.8000 ;
	    RECT 106.2000 63.8000 107.4000 64.1000 ;
	    RECT 107.8000 63.8000 108.2000 64.6000 ;
	    RECT 107.1000 63.5000 107.4000 63.8000 ;
	    RECT 107.1000 63.2000 108.9000 63.5000 ;
	    RECT 107.1000 63.1000 107.4000 63.2000 ;
	    RECT 107.0000 61.1000 107.4000 63.1000 ;
	    RECT 108.6000 63.1000 108.9000 63.2000 ;
	    RECT 108.6000 61.1000 109.0000 63.1000 ;
	    RECT 111.5000 61.1000 111.9000 64.8000 ;
	    RECT 112.3000 64.2000 112.6000 64.8000 ;
	    RECT 112.2000 63.8000 112.6000 64.2000 ;
	    RECT 113.5000 63.5000 113.8000 64.8000 ;
	    RECT 117.4000 64.7000 118.3000 65.1000 ;
	    RECT 119.0000 64.8000 119.4000 65.6000 ;
	    RECT 121.4000 65.2000 121.7000 66.8000 ;
	    RECT 123.0000 65.8000 123.4000 66.6000 ;
	    RECT 121.4000 64.8000 121.8000 65.2000 ;
	    RECT 123.7000 65.1000 124.0000 66.8000 ;
	    RECT 125.4000 66.1000 125.8000 69.9000 ;
	    RECT 127.0000 68.0000 127.4000 69.9000 ;
	    RECT 128.6000 68.0000 129.0000 69.9000 ;
	    RECT 127.0000 67.9000 129.0000 68.0000 ;
	    RECT 129.4000 67.9000 129.8000 69.9000 ;
	    RECT 130.3000 68.2000 130.7000 68.6000 ;
	    RECT 127.1000 67.7000 128.9000 67.9000 ;
	    RECT 126.2000 66.8000 126.6000 67.6000 ;
	    RECT 127.4000 67.2000 127.8000 67.4000 ;
	    RECT 129.4000 67.2000 129.7000 67.9000 ;
	    RECT 130.2000 67.8000 130.6000 68.2000 ;
	    RECT 131.0000 67.9000 131.4000 69.9000 ;
	    RECT 133.4000 67.9000 133.8000 69.9000 ;
	    RECT 134.2000 68.0000 134.6000 69.9000 ;
	    RECT 135.8000 68.0000 136.2000 69.9000 ;
	    RECT 134.2000 67.9000 136.2000 68.0000 ;
	    RECT 136.6000 68.0000 137.0000 69.9000 ;
	    RECT 138.2000 68.0000 138.6000 69.9000 ;
	    RECT 136.6000 67.9000 138.6000 68.0000 ;
	    RECT 139.0000 67.9000 139.4000 69.9000 ;
	    RECT 127.0000 66.9000 127.8000 67.2000 ;
	    RECT 127.0000 66.8000 127.4000 66.9000 ;
	    RECT 128.5000 66.8000 129.8000 67.2000 ;
	    RECT 126.2000 66.1000 126.6000 66.2000 ;
	    RECT 125.4000 65.8000 126.6000 66.1000 ;
	    RECT 127.8000 65.8000 128.2000 66.6000 ;
	    RECT 124.6000 65.1000 125.0000 65.2000 ;
	    RECT 123.5000 64.8000 124.0000 65.1000 ;
	    RECT 124.3000 64.8000 125.0000 65.1000 ;
	    RECT 114.2000 63.8000 114.6000 64.6000 ;
	    RECT 117.9000 64.1000 118.3000 64.7000 ;
	    RECT 120.6000 64.1000 121.0000 64.6000 ;
	    RECT 117.9000 63.8000 121.0000 64.1000 ;
	    RECT 113.5000 63.2000 115.3000 63.5000 ;
	    RECT 113.5000 63.1000 113.8000 63.2000 ;
	    RECT 113.4000 61.1000 113.8000 63.1000 ;
	    RECT 115.0000 63.1000 115.3000 63.2000 ;
	    RECT 115.0000 61.1000 115.4000 63.1000 ;
	    RECT 117.9000 61.1000 118.3000 63.8000 ;
	    RECT 121.4000 63.5000 121.7000 64.8000 ;
	    RECT 119.9000 63.2000 121.7000 63.5000 ;
	    RECT 119.8000 61.1000 120.2000 63.2000 ;
	    RECT 121.4000 63.1000 121.7000 63.2000 ;
	    RECT 121.4000 61.1000 121.8000 63.1000 ;
	    RECT 123.5000 61.1000 123.9000 64.8000 ;
	    RECT 124.3000 64.2000 124.6000 64.8000 ;
	    RECT 124.2000 63.8000 124.6000 64.2000 ;
	    RECT 125.4000 61.1000 125.8000 65.8000 ;
	    RECT 128.5000 65.1000 128.8000 66.8000 ;
	    RECT 130.2000 66.1000 130.6000 66.2000 ;
	    RECT 131.1000 66.1000 131.4000 67.9000 ;
	    RECT 133.5000 67.2000 133.8000 67.9000 ;
	    RECT 134.3000 67.7000 136.1000 67.9000 ;
	    RECT 136.7000 67.7000 138.5000 67.9000 ;
	    RECT 135.4000 67.2000 135.8000 67.4000 ;
	    RECT 137.0000 67.2000 137.4000 67.4000 ;
	    RECT 139.0000 67.2000 139.3000 67.9000 ;
	    RECT 131.8000 66.4000 132.2000 67.2000 ;
	    RECT 133.4000 66.8000 134.7000 67.2000 ;
	    RECT 135.4000 66.9000 136.2000 67.2000 ;
	    RECT 135.8000 66.8000 136.2000 66.9000 ;
	    RECT 136.6000 66.9000 137.4000 67.2000 ;
	    RECT 136.6000 66.8000 137.0000 66.9000 ;
	    RECT 138.1000 66.8000 139.4000 67.2000 ;
	    RECT 132.6000 66.1000 133.0000 66.2000 ;
	    RECT 130.2000 65.8000 131.4000 66.1000 ;
	    RECT 132.2000 65.8000 133.0000 66.1000 ;
	    RECT 129.4000 65.1000 129.8000 65.2000 ;
	    RECT 130.3000 65.1000 130.6000 65.8000 ;
	    RECT 132.2000 65.6000 132.6000 65.8000 ;
	    RECT 134.4000 65.2000 134.7000 66.8000 ;
	    RECT 135.0000 66.1000 135.4000 66.6000 ;
	    RECT 135.8000 66.1000 136.2000 66.2000 ;
	    RECT 135.0000 65.8000 136.2000 66.1000 ;
	    RECT 137.4000 65.8000 137.8000 66.6000 ;
	    RECT 133.4000 65.1000 133.8000 65.2000 ;
	    RECT 134.4000 65.1000 134.8000 65.2000 ;
	    RECT 138.1000 65.1000 138.4000 66.8000 ;
	    RECT 139.0000 65.1000 139.4000 65.2000 ;
	    RECT 128.3000 64.8000 128.8000 65.1000 ;
	    RECT 129.1000 64.8000 129.8000 65.1000 ;
	    RECT 128.3000 61.1000 128.7000 64.8000 ;
	    RECT 129.1000 64.2000 129.4000 64.8000 ;
	    RECT 129.0000 63.8000 129.4000 64.2000 ;
	    RECT 130.2000 61.1000 130.6000 65.1000 ;
	    RECT 131.0000 64.8000 133.0000 65.1000 ;
	    RECT 133.4000 64.8000 134.1000 65.1000 ;
	    RECT 134.4000 64.8000 134.9000 65.1000 ;
	    RECT 131.0000 61.1000 131.4000 64.8000 ;
	    RECT 132.6000 61.1000 133.0000 64.8000 ;
	    RECT 133.8000 64.2000 134.1000 64.8000 ;
	    RECT 133.4000 63.8000 134.2000 64.2000 ;
	    RECT 134.5000 61.1000 134.9000 64.8000 ;
	    RECT 137.9000 64.8000 138.4000 65.1000 ;
	    RECT 138.7000 64.8000 139.4000 65.1000 ;
	    RECT 137.9000 61.1000 138.3000 64.8000 ;
	    RECT 138.7000 64.2000 139.0000 64.8000 ;
	    RECT 138.6000 63.8000 139.0000 64.2000 ;
	    RECT 139.8000 61.1000 140.2000 69.9000 ;
	    RECT 142.7000 68.2000 143.1000 69.9000 ;
	    RECT 142.2000 67.9000 143.1000 68.2000 ;
	    RECT 140.6000 67.1000 141.0000 67.2000 ;
	    RECT 141.4000 67.1000 141.8000 67.6000 ;
	    RECT 140.6000 66.8000 141.8000 67.1000 ;
	    RECT 141.4000 65.8000 141.8000 66.2000 ;
	    RECT 141.4000 65.1000 141.7000 65.8000 ;
	    RECT 142.2000 65.1000 142.6000 67.9000 ;
	    RECT 141.4000 64.8000 142.6000 65.1000 ;
	    RECT 142.2000 61.1000 142.6000 64.8000 ;
	    RECT 143.8000 61.1000 144.2000 69.9000 ;
	    RECT 145.4000 67.6000 145.8000 69.9000 ;
	    RECT 145.4000 67.3000 146.5000 67.6000 ;
	    RECT 145.4000 65.8000 145.8000 66.6000 ;
	    RECT 146.2000 65.8000 146.5000 67.3000 ;
	    RECT 146.2000 65.4000 146.8000 65.8000 ;
	    RECT 146.2000 65.1000 146.5000 65.4000 ;
	    RECT 145.4000 64.8000 146.5000 65.1000 ;
	    RECT 145.4000 61.1000 145.8000 64.8000 ;
	    RECT 2.2000 56.2000 2.6000 59.9000 ;
	    RECT 4.6000 56.2000 5.0000 59.9000 ;
	    RECT 1.5000 55.9000 2.6000 56.2000 ;
	    RECT 3.9000 55.9000 5.0000 56.2000 ;
	    RECT 1.5000 55.6000 1.8000 55.9000 ;
	    RECT 3.9000 55.6000 4.2000 55.9000 ;
	    RECT 1.2000 55.2000 1.8000 55.6000 ;
	    RECT 3.6000 55.2000 4.2000 55.6000 ;
	    RECT 1.5000 53.7000 1.8000 55.2000 ;
	    RECT 2.2000 54.4000 2.6000 55.2000 ;
	    RECT 3.9000 53.7000 4.2000 55.2000 ;
	    RECT 4.6000 54.4000 5.0000 55.2000 ;
	    RECT 1.5000 53.4000 2.6000 53.7000 ;
	    RECT 3.9000 53.4000 5.0000 53.7000 ;
	    RECT 2.2000 51.1000 2.6000 53.4000 ;
	    RECT 4.6000 51.1000 5.0000 53.4000 ;
	    RECT 5.4000 52.4000 5.8000 53.2000 ;
	    RECT 6.2000 51.1000 6.6000 59.9000 ;
	    RECT 7.0000 55.9000 7.4000 59.9000 ;
	    RECT 8.6000 56.2000 9.0000 59.9000 ;
	    RECT 7.9000 55.9000 9.0000 56.2000 ;
	    RECT 7.0000 54.8000 7.3000 55.9000 ;
	    RECT 7.9000 55.6000 8.2000 55.9000 ;
	    RECT 7.6000 55.2000 8.2000 55.6000 ;
	    RECT 9.4000 55.6000 9.8000 59.9000 ;
	    RECT 11.5000 57.9000 12.1000 59.9000 ;
	    RECT 13.8000 57.9000 14.2000 59.9000 ;
	    RECT 16.0000 58.2000 16.4000 59.9000 ;
	    RECT 16.0000 57.9000 17.0000 58.2000 ;
	    RECT 11.8000 57.5000 12.2000 57.9000 ;
	    RECT 13.9000 57.6000 14.2000 57.9000 ;
	    RECT 13.5000 57.3000 15.3000 57.6000 ;
	    RECT 16.6000 57.5000 17.0000 57.9000 ;
	    RECT 13.5000 57.2000 13.9000 57.3000 ;
	    RECT 14.9000 57.2000 15.3000 57.3000 ;
	    RECT 11.0000 57.0000 11.7000 57.2000 ;
	    RECT 11.0000 56.8000 12.1000 57.0000 ;
	    RECT 11.4000 56.6000 12.1000 56.8000 ;
	    RECT 11.8000 56.1000 12.1000 56.6000 ;
	    RECT 12.9000 56.5000 14.0000 56.8000 ;
	    RECT 12.9000 56.4000 13.3000 56.5000 ;
	    RECT 11.8000 55.8000 13.0000 56.1000 ;
	    RECT 9.4000 55.3000 11.5000 55.6000 ;
	    RECT 7.0000 51.1000 7.4000 54.8000 ;
	    RECT 7.9000 53.7000 8.2000 55.2000 ;
	    RECT 8.6000 54.4000 9.0000 55.2000 ;
	    RECT 7.9000 53.4000 9.0000 53.7000 ;
	    RECT 8.6000 51.1000 9.0000 53.4000 ;
	    RECT 9.4000 53.6000 9.8000 55.3000 ;
	    RECT 11.1000 55.2000 11.5000 55.3000 ;
	    RECT 10.3000 54.9000 10.7000 55.0000 ;
	    RECT 10.3000 54.6000 12.2000 54.9000 ;
	    RECT 11.8000 54.5000 12.2000 54.6000 ;
	    RECT 12.7000 54.2000 13.0000 55.8000 ;
	    RECT 13.7000 55.9000 14.0000 56.5000 ;
	    RECT 14.3000 56.5000 14.7000 56.6000 ;
	    RECT 16.6000 56.5000 17.0000 56.6000 ;
	    RECT 14.3000 56.2000 17.0000 56.5000 ;
	    RECT 13.7000 55.7000 16.1000 55.9000 ;
	    RECT 18.2000 55.7000 18.6000 59.9000 ;
	    RECT 19.0000 56.2000 19.4000 59.9000 ;
	    RECT 19.9000 56.2000 20.3000 56.3000 ;
	    RECT 19.0000 55.9000 20.3000 56.2000 ;
	    RECT 21.2000 55.9000 22.0000 59.9000 ;
	    RECT 23.0000 56.2000 23.4000 56.3000 ;
	    RECT 23.8000 56.2000 24.2000 59.9000 ;
	    RECT 23.0000 55.9000 24.2000 56.2000 ;
	    RECT 13.7000 55.6000 18.6000 55.7000 ;
	    RECT 15.7000 55.5000 18.6000 55.6000 ;
	    RECT 15.8000 55.4000 18.6000 55.5000 ;
	    RECT 20.5000 55.2000 20.9000 55.3000 ;
	    RECT 21.5000 55.2000 21.8000 55.9000 ;
	    RECT 24.6000 55.7000 25.0000 59.9000 ;
	    RECT 26.8000 58.2000 27.2000 59.9000 ;
	    RECT 26.2000 57.9000 27.2000 58.2000 ;
	    RECT 29.0000 57.9000 29.4000 59.9000 ;
	    RECT 31.1000 57.9000 31.7000 59.9000 ;
	    RECT 26.2000 57.5000 26.6000 57.9000 ;
	    RECT 29.0000 57.6000 29.3000 57.9000 ;
	    RECT 27.9000 57.3000 29.7000 57.6000 ;
	    RECT 31.0000 57.5000 31.4000 57.9000 ;
	    RECT 27.9000 57.2000 28.3000 57.3000 ;
	    RECT 29.3000 57.2000 29.7000 57.3000 ;
	    RECT 26.2000 56.5000 26.6000 56.6000 ;
	    RECT 28.5000 56.5000 28.9000 56.6000 ;
	    RECT 26.2000 56.2000 28.9000 56.5000 ;
	    RECT 29.2000 56.5000 30.3000 56.8000 ;
	    RECT 29.2000 55.9000 29.5000 56.5000 ;
	    RECT 29.9000 56.4000 30.3000 56.5000 ;
	    RECT 31.1000 56.6000 31.8000 57.0000 ;
	    RECT 31.1000 56.1000 31.4000 56.6000 ;
	    RECT 27.1000 55.7000 29.5000 55.9000 ;
	    RECT 24.6000 55.6000 29.5000 55.7000 ;
	    RECT 30.2000 55.8000 31.4000 56.1000 ;
	    RECT 24.6000 55.5000 27.5000 55.6000 ;
	    RECT 24.6000 55.4000 27.4000 55.5000 ;
	    RECT 15.0000 55.1000 15.4000 55.2000 ;
	    RECT 15.0000 54.8000 17.5000 55.1000 ;
	    RECT 20.1000 54.9000 20.9000 55.2000 ;
	    RECT 21.4000 55.1000 21.8000 55.2000 ;
	    RECT 22.2000 55.1000 22.6000 55.2000 ;
	    RECT 27.8000 55.1000 28.2000 55.2000 ;
	    RECT 20.1000 54.8000 20.5000 54.9000 ;
	    RECT 21.4000 54.8000 22.6000 55.1000 ;
	    RECT 25.7000 54.8000 28.2000 55.1000 ;
	    RECT 15.8000 54.7000 16.2000 54.8000 ;
	    RECT 17.1000 54.7000 17.5000 54.8000 ;
	    RECT 20.8000 54.3000 21.2000 54.4000 ;
	    RECT 16.3000 54.2000 16.7000 54.3000 ;
	    RECT 19.8000 54.2000 21.2000 54.3000 ;
	    RECT 12.7000 53.9000 18.2000 54.2000 ;
	    RECT 12.9000 53.8000 13.3000 53.9000 ;
	    RECT 9.4000 53.3000 11.3000 53.6000 ;
	    RECT 9.4000 51.1000 9.8000 53.3000 ;
	    RECT 10.9000 53.2000 11.3000 53.3000 ;
	    RECT 15.8000 52.8000 16.1000 53.9000 ;
	    RECT 17.4000 53.8000 18.2000 53.9000 ;
	    RECT 19.0000 54.0000 21.2000 54.2000 ;
	    RECT 21.5000 54.2000 21.8000 54.8000 ;
	    RECT 25.7000 54.7000 26.1000 54.8000 ;
	    RECT 27.0000 54.7000 27.4000 54.8000 ;
	    RECT 26.5000 54.2000 26.9000 54.3000 ;
	    RECT 30.2000 54.2000 30.5000 55.8000 ;
	    RECT 33.4000 55.6000 33.8000 59.9000 ;
	    RECT 34.2000 56.2000 34.6000 59.9000 ;
	    RECT 34.2000 55.9000 35.3000 56.2000 ;
	    RECT 35.8000 55.9000 36.2000 59.9000 ;
	    RECT 37.4000 56.4000 37.8000 59.9000 ;
	    RECT 31.7000 55.3000 33.8000 55.6000 ;
	    RECT 31.7000 55.2000 32.1000 55.3000 ;
	    RECT 32.5000 54.9000 32.9000 55.0000 ;
	    RECT 31.0000 54.6000 32.9000 54.9000 ;
	    RECT 31.0000 54.5000 31.4000 54.6000 ;
	    RECT 19.0000 53.9000 20.1000 54.0000 ;
	    RECT 21.5000 53.9000 22.0000 54.2000 ;
	    RECT 19.0000 53.8000 19.8000 53.9000 ;
	    RECT 14.9000 52.7000 15.3000 52.8000 ;
	    RECT 11.8000 52.1000 12.2000 52.5000 ;
	    RECT 13.9000 52.4000 15.3000 52.7000 ;
	    RECT 15.8000 52.4000 16.2000 52.8000 ;
	    RECT 13.9000 52.1000 14.2000 52.4000 ;
	    RECT 16.6000 52.1000 17.0000 52.5000 ;
	    RECT 11.5000 51.8000 12.2000 52.1000 ;
	    RECT 11.5000 51.1000 12.1000 51.8000 ;
	    RECT 13.8000 51.1000 14.2000 52.1000 ;
	    RECT 16.0000 51.8000 17.0000 52.1000 ;
	    RECT 16.0000 51.1000 16.4000 51.8000 ;
	    RECT 18.2000 51.1000 18.6000 53.5000 ;
	    RECT 19.9000 53.4000 20.3000 53.5000 ;
	    RECT 19.0000 53.1000 20.3000 53.4000 ;
	    RECT 20.6000 53.2000 21.4000 53.6000 ;
	    RECT 19.0000 51.1000 19.4000 53.1000 ;
	    RECT 21.7000 52.9000 22.0000 53.9000 ;
	    RECT 22.4000 53.8000 22.8000 54.2000 ;
	    RECT 23.4000 53.8000 24.2000 54.2000 ;
	    RECT 25.0000 53.9000 30.5000 54.2000 ;
	    RECT 25.0000 53.8000 25.8000 53.9000 ;
	    RECT 22.4000 53.6000 22.7000 53.8000 ;
	    RECT 22.3000 53.2000 22.7000 53.6000 ;
	    RECT 23.0000 53.4000 23.4000 53.5000 ;
	    RECT 23.0000 53.1000 24.2000 53.4000 ;
	    RECT 21.2000 51.1000 22.0000 52.9000 ;
	    RECT 23.8000 51.1000 24.2000 53.1000 ;
	    RECT 24.6000 51.1000 25.0000 53.5000 ;
	    RECT 27.1000 52.8000 27.4000 53.9000 ;
	    RECT 29.9000 53.8000 30.3000 53.9000 ;
	    RECT 33.4000 53.6000 33.8000 55.3000 ;
	    RECT 35.0000 55.6000 35.3000 55.9000 ;
	    RECT 35.0000 55.2000 35.6000 55.6000 ;
	    RECT 34.2000 54.4000 34.6000 55.2000 ;
	    RECT 35.0000 53.7000 35.3000 55.2000 ;
	    RECT 35.9000 54.8000 36.2000 55.9000 ;
	    RECT 31.9000 53.3000 33.8000 53.6000 ;
	    RECT 31.9000 53.2000 32.3000 53.3000 ;
	    RECT 26.2000 52.1000 26.6000 52.5000 ;
	    RECT 27.0000 52.4000 27.4000 52.8000 ;
	    RECT 27.9000 52.7000 28.3000 52.8000 ;
	    RECT 27.9000 52.4000 29.3000 52.7000 ;
	    RECT 29.0000 52.1000 29.3000 52.4000 ;
	    RECT 31.0000 52.1000 31.4000 52.5000 ;
	    RECT 26.2000 51.8000 27.2000 52.1000 ;
	    RECT 26.8000 51.1000 27.2000 51.8000 ;
	    RECT 29.0000 51.1000 29.4000 52.1000 ;
	    RECT 31.0000 51.8000 31.7000 52.1000 ;
	    RECT 31.1000 51.1000 31.7000 51.8000 ;
	    RECT 33.4000 51.1000 33.8000 53.3000 ;
	    RECT 34.2000 53.4000 35.3000 53.7000 ;
	    RECT 34.2000 51.1000 34.6000 53.4000 ;
	    RECT 35.8000 51.1000 36.2000 54.8000 ;
	    RECT 37.3000 55.9000 37.8000 56.4000 ;
	    RECT 39.0000 56.2000 39.4000 59.9000 ;
	    RECT 38.1000 55.9000 39.4000 56.2000 ;
	    RECT 37.3000 54.2000 37.6000 55.9000 ;
	    RECT 38.1000 54.9000 38.4000 55.9000 ;
	    RECT 39.8000 55.8000 40.2000 56.6000 ;
	    RECT 37.9000 54.5000 38.4000 54.9000 ;
	    RECT 36.6000 54.1000 37.0000 54.2000 ;
	    RECT 37.3000 54.1000 37.8000 54.2000 ;
	    RECT 36.6000 53.8000 37.8000 54.1000 ;
	    RECT 37.3000 53.1000 37.6000 53.8000 ;
	    RECT 38.1000 53.7000 38.4000 54.5000 ;
	    RECT 38.9000 54.8000 39.4000 55.2000 ;
	    RECT 38.9000 54.4000 39.3000 54.8000 ;
	    RECT 38.1000 53.4000 39.4000 53.7000 ;
	    RECT 37.3000 52.8000 37.8000 53.1000 ;
	    RECT 37.4000 51.1000 37.8000 52.8000 ;
	    RECT 39.0000 51.1000 39.4000 53.4000 ;
	    RECT 40.6000 53.1000 41.0000 59.9000 ;
	    RECT 42.2000 56.2000 42.6000 59.9000 ;
	    RECT 43.0000 56.2000 43.4000 56.3000 ;
	    RECT 44.4000 56.2000 45.2000 59.9000 ;
	    RECT 42.2000 55.9000 43.4000 56.2000 ;
	    RECT 44.2000 55.9000 45.2000 56.2000 ;
	    RECT 46.3000 56.2000 46.7000 56.3000 ;
	    RECT 47.0000 56.2000 47.4000 59.9000 ;
	    RECT 46.3000 55.9000 47.4000 56.2000 ;
	    RECT 49.4000 56.2000 49.8000 59.9000 ;
	    RECT 50.1000 56.2000 50.5000 56.3000 ;
	    RECT 49.4000 55.9000 50.5000 56.2000 ;
	    RECT 51.6000 56.2000 52.4000 59.9000 ;
	    RECT 53.4000 56.2000 53.8000 56.3000 ;
	    RECT 54.2000 56.2000 54.6000 59.9000 ;
	    RECT 51.6000 55.9000 52.6000 56.2000 ;
	    RECT 53.4000 55.9000 54.6000 56.2000 ;
	    RECT 55.0000 56.2000 55.4000 59.9000 ;
	    RECT 56.6000 56.4000 57.0000 59.9000 ;
	    RECT 55.0000 55.9000 56.3000 56.2000 ;
	    RECT 56.6000 55.9000 57.1000 56.4000 ;
	    RECT 44.2000 55.2000 44.5000 55.9000 ;
	    RECT 46.3000 55.6000 46.6000 55.9000 ;
	    RECT 44.9000 55.3000 46.6000 55.6000 ;
	    RECT 50.2000 55.6000 50.5000 55.9000 ;
	    RECT 50.2000 55.3000 51.9000 55.6000 ;
	    RECT 44.9000 55.2000 45.3000 55.3000 ;
	    RECT 51.5000 55.2000 51.9000 55.3000 ;
	    RECT 52.3000 55.2000 52.6000 55.9000 ;
	    RECT 43.8000 54.9000 44.5000 55.2000 ;
	    RECT 46.0000 54.9000 46.4000 55.0000 ;
	    RECT 43.8000 54.8000 44.7000 54.9000 ;
	    RECT 44.2000 54.6000 44.7000 54.8000 ;
	    RECT 41.4000 53.4000 41.8000 54.2000 ;
	    RECT 42.2000 53.8000 43.0000 54.2000 ;
	    RECT 43.6000 53.8000 44.0000 54.2000 ;
	    RECT 43.7000 53.6000 44.0000 53.8000 ;
	    RECT 43.0000 53.4000 43.4000 53.5000 ;
	    RECT 40.1000 52.8000 41.0000 53.1000 ;
	    RECT 42.2000 53.1000 43.4000 53.4000 ;
	    RECT 43.7000 53.2000 44.1000 53.6000 ;
	    RECT 40.1000 51.1000 40.5000 52.8000 ;
	    RECT 42.2000 51.1000 42.6000 53.1000 ;
	    RECT 44.4000 52.9000 44.7000 54.6000 ;
	    RECT 45.1000 54.6000 46.4000 54.9000 ;
	    RECT 50.4000 54.9000 50.8000 55.0000 ;
	    RECT 52.3000 54.9000 53.0000 55.2000 ;
	    RECT 50.4000 54.6000 51.7000 54.9000 ;
	    RECT 45.1000 54.3000 45.4000 54.6000 ;
	    RECT 45.0000 53.9000 45.4000 54.3000 ;
	    RECT 51.4000 54.3000 51.7000 54.6000 ;
	    RECT 52.1000 54.8000 53.0000 54.9000 ;
	    RECT 54.2000 55.1000 54.6000 55.2000 ;
	    RECT 55.0000 55.1000 55.5000 55.2000 ;
	    RECT 54.2000 54.8000 55.5000 55.1000 ;
	    RECT 52.1000 54.6000 52.6000 54.8000 ;
	    RECT 46.6000 54.1000 47.4000 54.2000 ;
	    RECT 45.7000 53.8000 47.4000 54.1000 ;
	    RECT 49.4000 54.1000 50.2000 54.2000 ;
	    RECT 49.4000 53.8000 51.1000 54.1000 ;
	    RECT 51.4000 53.9000 51.8000 54.3000 ;
	    RECT 45.7000 53.6000 46.0000 53.8000 ;
	    RECT 45.0000 53.3000 46.0000 53.6000 ;
	    RECT 50.8000 53.6000 51.1000 53.8000 ;
	    RECT 46.3000 53.4000 46.7000 53.5000 ;
	    RECT 50.1000 53.4000 50.5000 53.5000 ;
	    RECT 45.0000 53.2000 45.8000 53.3000 ;
	    RECT 46.3000 53.1000 47.4000 53.4000 ;
	    RECT 44.4000 51.1000 45.2000 52.9000 ;
	    RECT 47.0000 51.1000 47.4000 53.1000 ;
	    RECT 49.4000 53.1000 50.5000 53.4000 ;
	    RECT 50.8000 53.3000 51.8000 53.6000 ;
	    RECT 51.0000 53.2000 51.8000 53.3000 ;
	    RECT 49.4000 51.1000 49.8000 53.1000 ;
	    RECT 52.1000 52.9000 52.4000 54.6000 ;
	    RECT 55.1000 54.4000 55.5000 54.8000 ;
	    RECT 56.0000 54.9000 56.3000 55.9000 ;
	    RECT 56.0000 54.5000 56.5000 54.9000 ;
	    RECT 52.8000 53.8000 53.2000 54.2000 ;
	    RECT 53.8000 53.8000 54.6000 54.2000 ;
	    RECT 52.8000 53.6000 53.1000 53.8000 ;
	    RECT 56.0000 53.7000 56.3000 54.5000 ;
	    RECT 56.8000 54.2000 57.1000 55.9000 ;
	    RECT 56.6000 53.8000 57.1000 54.2000 ;
	    RECT 52.7000 53.2000 53.1000 53.6000 ;
	    RECT 53.4000 53.4000 53.8000 53.5000 ;
	    RECT 55.0000 53.4000 56.3000 53.7000 ;
	    RECT 53.4000 53.1000 54.6000 53.4000 ;
	    RECT 51.6000 52.2000 52.4000 52.9000 ;
	    RECT 51.0000 51.8000 52.4000 52.2000 ;
	    RECT 51.6000 51.1000 52.4000 51.8000 ;
	    RECT 54.2000 51.1000 54.6000 53.1000 ;
	    RECT 55.0000 51.1000 55.4000 53.4000 ;
	    RECT 56.8000 53.1000 57.1000 53.8000 ;
	    RECT 56.6000 52.8000 57.1000 53.1000 ;
	    RECT 58.2000 55.8000 58.6000 59.9000 ;
	    RECT 59.8000 57.9000 60.2000 59.9000 ;
	    RECT 59.8000 55.8000 60.1000 57.9000 ;
	    RECT 62.7000 56.3000 63.1000 59.9000 ;
	    RECT 62.2000 55.9000 63.1000 56.3000 ;
	    RECT 63.8000 56.1000 64.2000 59.9000 ;
	    RECT 65.4000 56.1000 65.8000 56.6000 ;
	    RECT 58.2000 55.2000 58.5000 55.8000 ;
	    RECT 58.9000 55.5000 60.1000 55.8000 ;
	    RECT 58.2000 54.8000 58.6000 55.2000 ;
	    RECT 58.2000 53.1000 58.5000 54.8000 ;
	    RECT 58.9000 53.8000 59.2000 55.5000 ;
	    RECT 59.8000 54.8000 60.2000 55.2000 ;
	    RECT 59.8000 54.4000 60.1000 54.8000 ;
	    RECT 59.6000 54.0000 60.2000 54.4000 ;
	    RECT 60.6000 54.1000 61.0000 54.6000 ;
	    RECT 62.3000 54.2000 62.6000 55.9000 ;
	    RECT 63.8000 55.8000 65.8000 56.1000 ;
	    RECT 63.0000 54.8000 63.4000 55.6000 ;
	    RECT 62.2000 54.1000 62.6000 54.2000 ;
	    RECT 60.6000 53.8000 62.6000 54.1000 ;
	    RECT 58.8000 53.7000 59.2000 53.8000 ;
	    RECT 58.8000 53.5000 60.3000 53.7000 ;
	    RECT 58.8000 53.4000 60.9000 53.5000 ;
	    RECT 60.0000 53.2000 60.9000 53.4000 ;
	    RECT 60.6000 53.1000 60.9000 53.2000 ;
	    RECT 56.6000 51.1000 57.0000 52.8000 ;
	    RECT 58.2000 52.6000 58.9000 53.1000 ;
	    RECT 58.5000 51.1000 58.9000 52.6000 ;
	    RECT 60.6000 51.1000 61.0000 53.1000 ;
	    RECT 61.4000 52.4000 61.8000 53.2000 ;
	    RECT 62.3000 52.1000 62.6000 53.8000 ;
	    RECT 62.2000 51.1000 62.6000 52.1000 ;
	    RECT 63.8000 54.1000 64.2000 55.8000 ;
	    RECT 64.6000 54.1000 65.0000 54.2000 ;
	    RECT 63.8000 53.8000 65.0000 54.1000 ;
	    RECT 63.8000 51.1000 64.2000 53.8000 ;
	    RECT 64.6000 52.4000 65.0000 53.2000 ;
	    RECT 66.2000 53.1000 66.6000 59.9000 ;
	    RECT 68.6000 56.4000 69.0000 59.9000 ;
	    RECT 68.5000 55.9000 69.0000 56.4000 ;
	    RECT 70.2000 56.2000 70.6000 59.9000 ;
	    RECT 69.3000 55.9000 70.6000 56.2000 ;
	    RECT 68.5000 54.2000 68.8000 55.9000 ;
	    RECT 69.3000 54.9000 69.6000 55.9000 ;
	    RECT 69.1000 54.5000 69.6000 54.9000 ;
	    RECT 67.0000 53.4000 67.4000 54.2000 ;
	    RECT 67.8000 54.1000 68.2000 54.2000 ;
	    RECT 68.5000 54.1000 69.0000 54.2000 ;
	    RECT 67.8000 53.8000 69.0000 54.1000 ;
	    RECT 65.7000 52.8000 66.6000 53.1000 ;
	    RECT 68.5000 53.1000 68.8000 53.8000 ;
	    RECT 69.3000 53.7000 69.6000 54.5000 ;
	    RECT 70.1000 54.8000 70.6000 55.2000 ;
	    RECT 70.1000 54.4000 70.5000 54.8000 ;
	    RECT 69.3000 53.4000 70.6000 53.7000 ;
	    RECT 71.0000 53.4000 71.4000 54.2000 ;
	    RECT 68.5000 52.8000 69.0000 53.1000 ;
	    RECT 65.7000 51.1000 66.1000 52.8000 ;
	    RECT 68.6000 51.1000 69.0000 52.8000 ;
	    RECT 70.2000 51.1000 70.6000 53.4000 ;
	    RECT 71.8000 53.1000 72.2000 59.9000 ;
	    RECT 72.6000 55.8000 73.0000 56.6000 ;
	    RECT 74.7000 56.3000 75.1000 59.9000 ;
	    RECT 74.2000 55.9000 75.1000 56.3000 ;
	    RECT 76.1000 56.3000 76.5000 59.9000 ;
	    RECT 79.0000 56.4000 79.4000 59.9000 ;
	    RECT 76.1000 55.9000 77.0000 56.3000 ;
	    RECT 78.9000 55.9000 79.4000 56.4000 ;
	    RECT 80.6000 56.2000 81.0000 59.9000 ;
	    RECT 79.7000 55.9000 81.0000 56.2000 ;
	    RECT 82.7000 56.2000 83.1000 59.9000 ;
	    RECT 83.4000 56.8000 83.8000 57.2000 ;
	    RECT 83.5000 56.2000 83.8000 56.8000 ;
	    RECT 82.7000 55.9000 83.2000 56.2000 ;
	    RECT 83.5000 55.9000 84.2000 56.2000 ;
	    RECT 74.3000 54.2000 74.6000 55.9000 ;
	    RECT 75.0000 55.1000 75.4000 55.6000 ;
	    RECT 75.8000 55.1000 76.2000 55.6000 ;
	    RECT 75.0000 54.8000 76.2000 55.1000 ;
	    RECT 76.6000 54.2000 76.9000 55.9000 ;
	    RECT 78.9000 54.2000 79.2000 55.9000 ;
	    RECT 79.7000 54.9000 80.0000 55.9000 ;
	    RECT 79.5000 54.5000 80.0000 54.9000 ;
	    RECT 74.2000 54.1000 74.6000 54.2000 ;
	    RECT 75.0000 54.1000 75.4000 54.2000 ;
	    RECT 74.2000 53.8000 75.4000 54.1000 ;
	    RECT 76.6000 53.8000 77.0000 54.2000 ;
	    RECT 78.2000 54.1000 78.6000 54.2000 ;
	    RECT 78.9000 54.1000 79.4000 54.2000 ;
	    RECT 78.2000 53.8000 79.4000 54.1000 ;
	    RECT 73.4000 53.1000 73.8000 53.2000 ;
	    RECT 71.8000 52.8000 73.8000 53.1000 ;
	    RECT 72.3000 51.1000 72.7000 52.8000 ;
	    RECT 73.4000 52.4000 73.8000 52.8000 ;
	    RECT 74.3000 52.2000 74.6000 53.8000 ;
	    RECT 75.8000 53.1000 76.2000 53.2000 ;
	    RECT 76.6000 53.1000 76.9000 53.8000 ;
	    RECT 75.8000 52.8000 76.9000 53.1000 ;
	    RECT 74.2000 51.1000 74.6000 52.2000 ;
	    RECT 76.6000 52.1000 76.9000 52.8000 ;
	    RECT 77.4000 52.4000 77.8000 53.2000 ;
	    RECT 78.9000 53.1000 79.2000 53.8000 ;
	    RECT 79.7000 53.7000 80.0000 54.5000 ;
	    RECT 80.5000 54.8000 81.0000 55.2000 ;
	    RECT 81.4000 55.1000 81.8000 55.2000 ;
	    RECT 82.2000 55.1000 82.6000 55.2000 ;
	    RECT 81.4000 54.8000 82.6000 55.1000 ;
	    RECT 80.5000 54.4000 80.9000 54.8000 ;
	    RECT 82.2000 54.4000 82.6000 54.8000 ;
	    RECT 82.9000 54.2000 83.2000 55.9000 ;
	    RECT 83.8000 55.8000 84.2000 55.9000 ;
	    RECT 84.6000 55.8000 85.0000 56.6000 ;
	    RECT 83.8000 55.1000 84.1000 55.8000 ;
	    RECT 85.4000 55.1000 85.8000 59.9000 ;
	    RECT 83.8000 54.8000 85.8000 55.1000 ;
	    RECT 81.4000 54.1000 81.8000 54.2000 ;
	    RECT 81.4000 53.8000 82.2000 54.1000 ;
	    RECT 82.9000 53.8000 84.2000 54.2000 ;
	    RECT 79.7000 53.4000 81.0000 53.7000 ;
	    RECT 81.8000 53.6000 82.2000 53.8000 ;
	    RECT 78.9000 52.8000 79.4000 53.1000 ;
	    RECT 76.6000 51.1000 77.0000 52.1000 ;
	    RECT 79.0000 51.1000 79.4000 52.8000 ;
	    RECT 80.6000 51.1000 81.0000 53.4000 ;
	    RECT 81.5000 53.1000 83.3000 53.3000 ;
	    RECT 83.8000 53.1000 84.1000 53.8000 ;
	    RECT 85.4000 53.1000 85.8000 54.8000 ;
	    RECT 87.8000 55.1000 88.2000 59.9000 ;
	    RECT 88.9000 56.3000 89.3000 59.9000 ;
	    RECT 91.0000 59.6000 93.0000 59.9000 ;
	    RECT 88.9000 55.9000 89.8000 56.3000 ;
	    RECT 91.0000 55.9000 91.4000 59.6000 ;
	    RECT 91.8000 55.9000 92.2000 59.3000 ;
	    RECT 92.6000 56.2000 93.0000 59.6000 ;
	    RECT 94.2000 56.2000 94.6000 59.9000 ;
	    RECT 92.6000 55.9000 94.6000 56.2000 ;
	    RECT 88.6000 55.1000 89.0000 55.6000 ;
	    RECT 87.8000 54.8000 89.0000 55.1000 ;
	    RECT 86.2000 54.1000 86.6000 54.2000 ;
	    RECT 87.0000 54.1000 87.4000 54.2000 ;
	    RECT 86.2000 53.8000 87.4000 54.1000 ;
	    RECT 86.2000 53.4000 86.6000 53.8000 ;
	    RECT 81.4000 53.0000 83.4000 53.1000 ;
	    RECT 81.4000 51.1000 81.8000 53.0000 ;
	    RECT 83.0000 51.1000 83.4000 53.0000 ;
	    RECT 83.8000 51.1000 84.2000 53.1000 ;
	    RECT 84.9000 52.8000 85.8000 53.1000 ;
	    RECT 84.9000 51.1000 85.3000 52.8000 ;
	    RECT 87.0000 52.4000 87.4000 53.2000 ;
	    RECT 87.8000 51.1000 88.2000 54.8000 ;
	    RECT 89.4000 54.2000 89.7000 55.9000 ;
	    RECT 91.9000 55.6000 92.2000 55.9000 ;
	    RECT 96.6000 55.6000 97.0000 59.9000 ;
	    RECT 98.7000 57.9000 99.3000 59.9000 ;
	    RECT 101.0000 57.9000 101.4000 59.9000 ;
	    RECT 103.2000 58.2000 103.6000 59.9000 ;
	    RECT 103.2000 57.9000 104.2000 58.2000 ;
	    RECT 99.0000 57.5000 99.4000 57.9000 ;
	    RECT 101.1000 57.6000 101.4000 57.9000 ;
	    RECT 100.7000 57.3000 102.5000 57.6000 ;
	    RECT 103.8000 57.5000 104.2000 57.9000 ;
	    RECT 100.7000 57.2000 101.1000 57.3000 ;
	    RECT 102.1000 57.2000 102.5000 57.3000 ;
	    RECT 98.6000 56.6000 99.3000 57.0000 ;
	    RECT 99.0000 56.1000 99.3000 56.6000 ;
	    RECT 100.1000 56.5000 101.2000 56.8000 ;
	    RECT 100.1000 56.4000 100.5000 56.5000 ;
	    RECT 99.0000 55.8000 100.2000 56.1000 ;
	    RECT 91.0000 54.8000 91.4000 55.6000 ;
	    RECT 91.9000 55.3000 92.9000 55.6000 ;
	    RECT 92.6000 55.2000 92.9000 55.3000 ;
	    RECT 93.8000 55.2000 94.2000 55.4000 ;
	    RECT 96.6000 55.3000 98.7000 55.6000 ;
	    RECT 92.6000 54.8000 93.0000 55.2000 ;
	    RECT 93.8000 54.9000 94.6000 55.2000 ;
	    RECT 94.2000 54.8000 94.6000 54.9000 ;
	    RECT 91.9000 54.4000 92.3000 54.8000 ;
	    RECT 91.9000 54.2000 92.2000 54.4000 ;
	    RECT 89.4000 53.8000 89.8000 54.2000 ;
	    RECT 91.8000 53.8000 92.2000 54.2000 ;
	    RECT 89.4000 52.2000 89.7000 53.8000 ;
	    RECT 90.2000 52.4000 90.6000 53.2000 ;
	    RECT 92.6000 53.1000 92.9000 54.8000 ;
	    RECT 93.4000 53.8000 93.8000 54.6000 ;
	    RECT 96.6000 53.6000 97.0000 55.3000 ;
	    RECT 98.3000 55.2000 98.7000 55.3000 ;
	    RECT 97.5000 54.9000 97.9000 55.0000 ;
	    RECT 97.5000 54.6000 99.4000 54.9000 ;
	    RECT 99.0000 54.5000 99.4000 54.6000 ;
	    RECT 99.9000 54.2000 100.2000 55.8000 ;
	    RECT 100.9000 55.9000 101.2000 56.5000 ;
	    RECT 101.5000 56.5000 101.9000 56.6000 ;
	    RECT 103.8000 56.5000 104.2000 56.6000 ;
	    RECT 101.5000 56.2000 104.2000 56.5000 ;
	    RECT 100.9000 55.7000 103.3000 55.9000 ;
	    RECT 105.4000 55.7000 105.8000 59.9000 ;
	    RECT 106.5000 56.3000 106.9000 59.9000 ;
	    RECT 106.5000 55.9000 107.4000 56.3000 ;
	    RECT 108.6000 56.2000 109.0000 59.9000 ;
	    RECT 110.2000 56.4000 110.6000 59.9000 ;
	    RECT 112.9000 57.2000 113.3000 59.9000 ;
	    RECT 115.8000 57.9000 116.2000 59.9000 ;
	    RECT 112.2000 56.8000 112.6000 57.2000 ;
	    RECT 112.9000 56.8000 113.8000 57.2000 ;
	    RECT 108.6000 55.9000 109.9000 56.2000 ;
	    RECT 110.2000 55.9000 110.7000 56.4000 ;
	    RECT 112.2000 56.2000 112.5000 56.8000 ;
	    RECT 112.9000 56.2000 113.3000 56.8000 ;
	    RECT 100.9000 55.6000 105.8000 55.7000 ;
	    RECT 102.9000 55.5000 105.8000 55.6000 ;
	    RECT 103.0000 55.4000 105.8000 55.5000 ;
	    RECT 102.2000 55.1000 102.6000 55.2000 ;
	    RECT 102.2000 54.8000 104.7000 55.1000 ;
	    RECT 106.2000 54.8000 106.6000 55.6000 ;
	    RECT 103.0000 54.7000 103.4000 54.8000 ;
	    RECT 104.3000 54.7000 104.7000 54.8000 ;
	    RECT 103.5000 54.2000 103.9000 54.3000 ;
	    RECT 107.0000 54.2000 107.3000 55.9000 ;
	    RECT 108.6000 54.8000 109.1000 55.2000 ;
	    RECT 108.7000 54.4000 109.1000 54.8000 ;
	    RECT 109.6000 54.9000 109.9000 55.9000 ;
	    RECT 109.6000 54.5000 110.1000 54.9000 ;
	    RECT 99.9000 53.9000 105.4000 54.2000 ;
	    RECT 100.1000 53.8000 100.5000 53.9000 ;
	    RECT 96.6000 53.3000 98.5000 53.6000 ;
	    RECT 89.4000 51.1000 89.8000 52.2000 ;
	    RECT 92.3000 51.1000 93.1000 53.1000 ;
	    RECT 96.6000 51.1000 97.0000 53.3000 ;
	    RECT 98.1000 53.2000 98.5000 53.3000 ;
	    RECT 103.0000 52.8000 103.3000 53.9000 ;
	    RECT 104.6000 53.8000 105.4000 53.9000 ;
	    RECT 107.0000 53.8000 107.4000 54.2000 ;
	    RECT 102.1000 52.7000 102.5000 52.8000 ;
	    RECT 99.0000 52.1000 99.4000 52.5000 ;
	    RECT 101.1000 52.4000 102.5000 52.7000 ;
	    RECT 103.0000 52.4000 103.4000 52.8000 ;
	    RECT 101.1000 52.1000 101.4000 52.4000 ;
	    RECT 103.8000 52.1000 104.2000 52.5000 ;
	    RECT 98.7000 51.8000 99.4000 52.1000 ;
	    RECT 98.7000 51.1000 99.3000 51.8000 ;
	    RECT 101.0000 51.1000 101.4000 52.1000 ;
	    RECT 103.2000 51.8000 104.2000 52.1000 ;
	    RECT 103.2000 51.1000 103.6000 51.8000 ;
	    RECT 105.4000 51.1000 105.8000 53.5000 ;
	    RECT 107.0000 52.2000 107.3000 53.8000 ;
	    RECT 109.6000 53.7000 109.9000 54.5000 ;
	    RECT 110.4000 54.2000 110.7000 55.9000 ;
	    RECT 111.8000 55.9000 112.5000 56.2000 ;
	    RECT 112.8000 55.9000 113.3000 56.2000 ;
	    RECT 111.8000 55.8000 112.2000 55.9000 ;
	    RECT 112.8000 54.2000 113.1000 55.9000 ;
	    RECT 115.9000 55.8000 116.2000 57.9000 ;
	    RECT 117.4000 55.9000 117.8000 59.9000 ;
	    RECT 119.5000 59.2000 119.9000 59.9000 ;
	    RECT 119.0000 58.8000 119.9000 59.2000 ;
	    RECT 119.5000 56.2000 119.9000 58.8000 ;
	    RECT 120.2000 56.8000 120.6000 57.2000 ;
	    RECT 120.3000 56.2000 120.6000 56.8000 ;
	    RECT 121.8000 56.8000 122.2000 57.2000 ;
	    RECT 121.8000 56.2000 122.1000 56.8000 ;
	    RECT 122.5000 56.2000 122.9000 59.9000 ;
	    RECT 125.9000 57.2000 126.3000 59.9000 ;
	    RECT 125.4000 56.8000 126.3000 57.2000 ;
	    RECT 126.6000 56.8000 127.0000 57.2000 ;
	    RECT 119.5000 55.9000 120.0000 56.2000 ;
	    RECT 120.3000 55.9000 121.0000 56.2000 ;
	    RECT 115.9000 55.5000 117.1000 55.8000 ;
	    RECT 113.4000 54.4000 113.8000 55.2000 ;
	    RECT 115.8000 54.8000 116.2000 55.2000 ;
	    RECT 110.2000 53.8000 110.7000 54.2000 ;
	    RECT 111.8000 53.8000 113.1000 54.2000 ;
	    RECT 114.2000 54.1000 114.6000 54.2000 ;
	    RECT 115.0000 54.1000 115.4000 54.6000 ;
	    RECT 115.9000 54.4000 116.2000 54.8000 ;
	    RECT 115.9000 54.1000 116.4000 54.4000 ;
	    RECT 113.8000 53.8000 115.4000 54.1000 ;
	    RECT 116.0000 54.0000 116.4000 54.1000 ;
	    RECT 116.8000 53.8000 117.1000 55.5000 ;
	    RECT 117.5000 55.2000 117.8000 55.9000 ;
	    RECT 117.4000 55.1000 117.8000 55.2000 ;
	    RECT 117.4000 54.8000 118.5000 55.1000 ;
	    RECT 108.6000 53.4000 109.9000 53.7000 ;
	    RECT 107.8000 52.4000 108.2000 53.2000 ;
	    RECT 107.0000 51.1000 107.4000 52.2000 ;
	    RECT 108.6000 51.1000 109.0000 53.4000 ;
	    RECT 110.4000 53.1000 110.7000 53.8000 ;
	    RECT 111.9000 53.1000 112.2000 53.8000 ;
	    RECT 113.8000 53.6000 114.2000 53.8000 ;
	    RECT 116.8000 53.7000 117.2000 53.8000 ;
	    RECT 115.7000 53.5000 117.2000 53.7000 ;
	    RECT 115.1000 53.4000 117.2000 53.5000 ;
	    RECT 112.7000 53.1000 114.5000 53.3000 ;
	    RECT 115.1000 53.2000 116.0000 53.4000 ;
	    RECT 115.1000 53.1000 115.4000 53.2000 ;
	    RECT 117.5000 53.1000 117.8000 54.8000 ;
	    RECT 118.2000 54.2000 118.5000 54.8000 ;
	    RECT 119.0000 54.4000 119.4000 55.2000 ;
	    RECT 119.7000 54.2000 120.0000 55.9000 ;
	    RECT 120.6000 55.8000 121.0000 55.9000 ;
	    RECT 121.4000 55.9000 122.1000 56.2000 ;
	    RECT 122.4000 55.9000 122.9000 56.2000 ;
	    RECT 125.9000 56.2000 126.3000 56.8000 ;
	    RECT 126.7000 56.2000 127.0000 56.8000 ;
	    RECT 125.9000 55.9000 126.4000 56.2000 ;
	    RECT 126.7000 56.1000 127.4000 56.2000 ;
	    RECT 128.6000 56.1000 129.0000 59.9000 ;
	    RECT 126.7000 55.9000 129.0000 56.1000 ;
	    RECT 130.2000 56.2000 130.6000 59.9000 ;
	    RECT 131.8000 56.2000 132.2000 59.9000 ;
	    RECT 130.2000 55.9000 132.2000 56.2000 ;
	    RECT 132.6000 55.9000 133.0000 59.9000 ;
	    RECT 133.4000 55.9000 133.8000 59.9000 ;
	    RECT 134.2000 56.2000 134.6000 59.9000 ;
	    RECT 135.8000 56.2000 136.2000 59.9000 ;
	    RECT 134.2000 55.9000 136.2000 56.2000 ;
	    RECT 121.4000 55.8000 121.8000 55.9000 ;
	    RECT 120.6000 55.1000 120.9000 55.8000 ;
	    RECT 122.4000 55.1000 122.7000 55.9000 ;
	    RECT 120.6000 54.8000 122.7000 55.1000 ;
	    RECT 122.4000 54.2000 122.7000 54.8000 ;
	    RECT 123.0000 55.1000 123.4000 55.2000 ;
	    RECT 123.8000 55.1000 124.2000 55.2000 ;
	    RECT 123.0000 54.8000 124.2000 55.1000 ;
	    RECT 123.0000 54.4000 123.4000 54.8000 ;
	    RECT 125.4000 54.4000 125.8000 55.2000 ;
	    RECT 126.1000 54.2000 126.4000 55.9000 ;
	    RECT 127.0000 55.8000 129.0000 55.9000 ;
	    RECT 118.2000 54.1000 118.6000 54.2000 ;
	    RECT 118.2000 53.8000 119.0000 54.1000 ;
	    RECT 119.7000 53.8000 121.0000 54.2000 ;
	    RECT 121.4000 53.8000 122.7000 54.2000 ;
	    RECT 123.8000 54.1000 124.2000 54.2000 ;
	    RECT 123.4000 53.8000 124.2000 54.1000 ;
	    RECT 124.6000 54.1000 125.0000 54.2000 ;
	    RECT 124.6000 53.8000 125.4000 54.1000 ;
	    RECT 126.1000 53.8000 127.4000 54.2000 ;
	    RECT 118.6000 53.6000 119.0000 53.8000 ;
	    RECT 118.3000 53.1000 120.1000 53.3000 ;
	    RECT 120.6000 53.1000 120.9000 53.8000 ;
	    RECT 121.5000 53.1000 121.8000 53.8000 ;
	    RECT 123.4000 53.6000 123.8000 53.8000 ;
	    RECT 125.0000 53.6000 125.4000 53.8000 ;
	    RECT 122.3000 53.1000 124.1000 53.3000 ;
	    RECT 124.7000 53.1000 126.5000 53.3000 ;
	    RECT 127.0000 53.1000 127.3000 53.8000 ;
	    RECT 127.8000 53.4000 128.2000 54.2000 ;
	    RECT 128.6000 53.1000 129.0000 55.8000 ;
	    RECT 130.6000 55.2000 131.0000 55.4000 ;
	    RECT 132.6000 55.2000 132.9000 55.9000 ;
	    RECT 133.5000 55.2000 133.8000 55.9000 ;
	    RECT 135.4000 55.2000 135.8000 55.4000 ;
	    RECT 130.2000 54.9000 131.0000 55.2000 ;
	    RECT 131.8000 54.9000 133.0000 55.2000 ;
	    RECT 130.2000 54.8000 130.6000 54.9000 ;
	    RECT 131.0000 53.8000 131.4000 54.6000 ;
	    RECT 131.8000 53.1000 132.1000 54.9000 ;
	    RECT 132.6000 54.8000 133.0000 54.9000 ;
	    RECT 133.4000 54.9000 134.6000 55.2000 ;
	    RECT 135.4000 54.9000 136.2000 55.2000 ;
	    RECT 133.4000 54.8000 133.8000 54.9000 ;
	    RECT 132.6000 53.1000 133.0000 53.2000 ;
	    RECT 133.4000 53.1000 133.8000 53.2000 ;
	    RECT 134.3000 53.1000 134.6000 54.9000 ;
	    RECT 135.8000 54.8000 136.2000 54.9000 ;
	    RECT 135.0000 54.1000 135.4000 54.6000 ;
	    RECT 136.6000 54.1000 137.0000 59.9000 ;
	    RECT 138.2000 56.2000 138.6000 59.9000 ;
	    RECT 138.2000 55.9000 139.3000 56.2000 ;
	    RECT 139.0000 55.6000 139.3000 55.9000 ;
	    RECT 139.0000 55.2000 139.6000 55.6000 ;
	    RECT 137.4000 55.1000 137.8000 55.2000 ;
	    RECT 138.2000 55.1000 138.6000 55.2000 ;
	    RECT 137.4000 54.8000 138.6000 55.1000 ;
	    RECT 138.2000 54.4000 138.6000 54.8000 ;
	    RECT 135.0000 53.8000 137.0000 54.1000 ;
	    RECT 110.2000 52.8000 110.7000 53.1000 ;
	    RECT 110.2000 51.1000 110.6000 52.8000 ;
	    RECT 111.8000 51.1000 112.2000 53.1000 ;
	    RECT 112.6000 53.0000 114.6000 53.1000 ;
	    RECT 112.6000 51.1000 113.0000 53.0000 ;
	    RECT 114.2000 51.1000 114.6000 53.0000 ;
	    RECT 115.0000 51.1000 115.4000 53.1000 ;
	    RECT 117.1000 52.6000 117.8000 53.1000 ;
	    RECT 118.2000 53.0000 120.2000 53.1000 ;
	    RECT 117.1000 51.1000 117.5000 52.6000 ;
	    RECT 118.2000 51.1000 118.6000 53.0000 ;
	    RECT 119.8000 51.1000 120.2000 53.0000 ;
	    RECT 120.6000 51.1000 121.0000 53.1000 ;
	    RECT 121.4000 51.1000 121.8000 53.1000 ;
	    RECT 122.2000 53.0000 124.2000 53.1000 ;
	    RECT 122.2000 51.1000 122.6000 53.0000 ;
	    RECT 123.8000 51.1000 124.2000 53.0000 ;
	    RECT 124.6000 53.0000 126.6000 53.1000 ;
	    RECT 124.6000 51.1000 125.0000 53.0000 ;
	    RECT 126.2000 51.1000 126.6000 53.0000 ;
	    RECT 127.0000 51.1000 127.4000 53.1000 ;
	    RECT 128.6000 52.8000 129.5000 53.1000 ;
	    RECT 129.1000 51.1000 129.5000 52.8000 ;
	    RECT 131.8000 51.1000 132.2000 53.1000 ;
	    RECT 132.6000 52.8000 133.8000 53.1000 ;
	    RECT 132.5000 52.4000 132.9000 52.8000 ;
	    RECT 133.5000 52.4000 133.9000 52.8000 ;
	    RECT 134.2000 51.1000 134.6000 53.1000 ;
	    RECT 136.6000 51.1000 137.0000 53.8000 ;
	    RECT 139.0000 53.7000 139.3000 55.2000 ;
	    RECT 138.2000 53.4000 139.3000 53.7000 ;
	    RECT 140.6000 53.4000 141.0000 54.2000 ;
	    RECT 138.2000 51.1000 138.6000 53.4000 ;
	    RECT 141.4000 53.1000 141.8000 59.9000 ;
	    RECT 143.0000 56.2000 143.4000 59.9000 ;
	    RECT 143.0000 55.9000 144.1000 56.2000 ;
	    RECT 143.8000 55.6000 144.1000 55.9000 ;
	    RECT 143.8000 55.2000 144.4000 55.6000 ;
	    RECT 142.2000 55.1000 142.6000 55.2000 ;
	    RECT 143.0000 55.1000 143.4000 55.2000 ;
	    RECT 142.2000 54.8000 143.4000 55.1000 ;
	    RECT 143.0000 54.4000 143.4000 54.8000 ;
	    RECT 143.8000 53.7000 144.1000 55.2000 ;
	    RECT 143.0000 53.4000 144.1000 53.7000 ;
	    RECT 145.4000 53.4000 145.8000 54.2000 ;
	    RECT 141.4000 52.8000 142.3000 53.1000 ;
	    RECT 141.9000 52.2000 142.3000 52.8000 ;
	    RECT 141.4000 51.8000 142.3000 52.2000 ;
	    RECT 141.9000 51.1000 142.3000 51.8000 ;
	    RECT 143.0000 51.1000 143.4000 53.4000 ;
	    RECT 146.2000 53.1000 146.6000 59.9000 ;
	    RECT 146.2000 52.8000 147.1000 53.1000 ;
	    RECT 146.7000 51.1000 147.1000 52.8000 ;
	    RECT 0.6000 47.7000 1.0000 49.9000 ;
	    RECT 2.7000 49.2000 3.3000 49.9000 ;
	    RECT 2.7000 48.9000 3.4000 49.2000 ;
	    RECT 5.0000 48.9000 5.4000 49.9000 ;
	    RECT 7.2000 49.2000 7.6000 49.9000 ;
	    RECT 7.2000 48.9000 8.2000 49.2000 ;
	    RECT 3.0000 48.5000 3.4000 48.9000 ;
	    RECT 5.1000 48.6000 5.4000 48.9000 ;
	    RECT 5.1000 48.3000 6.5000 48.6000 ;
	    RECT 6.1000 48.2000 6.5000 48.3000 ;
	    RECT 7.0000 48.2000 7.4000 48.6000 ;
	    RECT 7.8000 48.5000 8.2000 48.9000 ;
	    RECT 2.1000 47.7000 2.5000 47.8000 ;
	    RECT 0.6000 47.4000 2.5000 47.7000 ;
	    RECT 0.6000 45.7000 1.0000 47.4000 ;
	    RECT 4.1000 47.1000 4.5000 47.2000 ;
	    RECT 7.0000 47.1000 7.3000 48.2000 ;
	    RECT 9.4000 47.5000 9.8000 49.9000 ;
	    RECT 11.0000 48.9000 11.4000 49.9000 ;
	    RECT 10.2000 47.8000 10.6000 48.6000 ;
	    RECT 11.1000 47.2000 11.4000 48.9000 ;
	    RECT 12.6000 47.6000 13.0000 49.9000 ;
	    RECT 12.6000 47.3000 13.7000 47.6000 ;
	    RECT 8.6000 47.1000 9.4000 47.2000 ;
	    RECT 11.0000 47.1000 11.4000 47.2000 ;
	    RECT 3.9000 46.8000 9.4000 47.1000 ;
	    RECT 10.2000 46.8000 11.4000 47.1000 ;
	    RECT 3.0000 46.4000 3.4000 46.5000 ;
	    RECT 1.5000 46.1000 3.4000 46.4000 ;
	    RECT 1.5000 46.0000 1.9000 46.1000 ;
	    RECT 2.3000 45.7000 2.7000 45.8000 ;
	    RECT 0.6000 45.4000 2.7000 45.7000 ;
	    RECT 0.6000 41.1000 1.0000 45.4000 ;
	    RECT 3.9000 45.2000 4.2000 46.8000 ;
	    RECT 7.5000 46.7000 7.9000 46.8000 ;
	    RECT 7.0000 46.2000 7.4000 46.3000 ;
	    RECT 8.3000 46.2000 8.7000 46.3000 ;
	    RECT 6.2000 45.9000 8.7000 46.2000 ;
	    RECT 10.2000 46.2000 10.5000 46.8000 ;
	    RECT 6.2000 45.8000 6.6000 45.9000 ;
	    RECT 10.2000 45.8000 10.6000 46.2000 ;
	    RECT 7.0000 45.5000 9.8000 45.6000 ;
	    RECT 6.9000 45.4000 9.8000 45.5000 ;
	    RECT 3.0000 44.9000 4.2000 45.2000 ;
	    RECT 4.9000 45.3000 9.8000 45.4000 ;
	    RECT 4.9000 45.1000 7.3000 45.3000 ;
	    RECT 3.0000 44.4000 3.3000 44.9000 ;
	    RECT 2.6000 44.0000 3.3000 44.4000 ;
	    RECT 4.1000 44.5000 4.5000 44.6000 ;
	    RECT 4.9000 44.5000 5.2000 45.1000 ;
	    RECT 4.1000 44.2000 5.2000 44.5000 ;
	    RECT 5.5000 44.5000 8.2000 44.8000 ;
	    RECT 5.5000 44.4000 5.9000 44.5000 ;
	    RECT 7.8000 44.4000 8.2000 44.5000 ;
	    RECT 4.7000 43.7000 5.1000 43.8000 ;
	    RECT 6.1000 43.7000 6.5000 43.8000 ;
	    RECT 3.0000 43.1000 3.4000 43.5000 ;
	    RECT 4.7000 43.4000 6.5000 43.7000 ;
	    RECT 5.1000 43.1000 5.4000 43.4000 ;
	    RECT 7.8000 43.1000 8.2000 43.5000 ;
	    RECT 2.7000 41.1000 3.3000 43.1000 ;
	    RECT 5.0000 41.1000 5.4000 43.1000 ;
	    RECT 7.2000 42.8000 8.2000 43.1000 ;
	    RECT 7.2000 41.1000 7.6000 42.8000 ;
	    RECT 9.4000 41.1000 9.8000 45.3000 ;
	    RECT 11.1000 45.1000 11.4000 46.8000 ;
	    RECT 11.8000 45.4000 12.2000 46.2000 ;
	    RECT 12.6000 45.8000 13.0000 46.6000 ;
	    RECT 13.4000 45.8000 13.7000 47.3000 ;
	    RECT 14.2000 46.2000 14.6000 49.9000 ;
	    RECT 13.4000 45.4000 14.0000 45.8000 ;
	    RECT 13.4000 45.1000 13.7000 45.4000 ;
	    RECT 14.3000 45.1000 14.6000 46.2000 ;
	    RECT 11.0000 44.7000 11.9000 45.1000 ;
	    RECT 11.5000 41.1000 11.9000 44.7000 ;
	    RECT 12.6000 44.8000 13.7000 45.1000 ;
	    RECT 12.6000 41.1000 13.0000 44.8000 ;
	    RECT 14.2000 41.1000 14.6000 45.1000 ;
	    RECT 15.0000 46.2000 15.4000 49.9000 ;
	    RECT 16.6000 47.6000 17.0000 49.9000 ;
	    RECT 18.2000 48.2000 18.6000 49.9000 ;
	    RECT 15.9000 47.3000 17.0000 47.6000 ;
	    RECT 18.1000 47.9000 18.6000 48.2000 ;
	    RECT 15.0000 45.1000 15.3000 46.2000 ;
	    RECT 15.9000 45.8000 16.2000 47.3000 ;
	    RECT 18.1000 47.2000 18.4000 47.9000 ;
	    RECT 19.8000 47.6000 20.2000 49.9000 ;
	    RECT 18.9000 47.3000 20.2000 47.6000 ;
	    RECT 20.6000 47.6000 21.0000 49.9000 ;
	    RECT 20.6000 47.3000 21.7000 47.6000 ;
	    RECT 17.4000 47.1000 17.8000 47.2000 ;
	    RECT 18.1000 47.1000 18.6000 47.2000 ;
	    RECT 17.4000 46.8000 18.6000 47.1000 ;
	    RECT 16.6000 45.8000 17.0000 46.6000 ;
	    RECT 15.6000 45.4000 16.2000 45.8000 ;
	    RECT 15.9000 45.1000 16.2000 45.4000 ;
	    RECT 18.1000 45.1000 18.4000 46.8000 ;
	    RECT 18.9000 46.5000 19.2000 47.3000 ;
	    RECT 18.7000 46.1000 19.2000 46.5000 ;
	    RECT 18.9000 45.1000 19.2000 46.1000 ;
	    RECT 20.6000 45.8000 21.0000 46.6000 ;
	    RECT 21.4000 45.8000 21.7000 47.3000 ;
	    RECT 22.2000 46.2000 22.6000 49.9000 ;
	    RECT 21.4000 45.4000 22.0000 45.8000 ;
	    RECT 21.4000 45.1000 21.7000 45.4000 ;
	    RECT 22.3000 45.1000 22.6000 46.2000 ;
	    RECT 15.0000 41.1000 15.4000 45.1000 ;
	    RECT 15.9000 44.8000 17.0000 45.1000 ;
	    RECT 16.6000 41.1000 17.0000 44.8000 ;
	    RECT 18.1000 44.6000 18.6000 45.1000 ;
	    RECT 18.9000 44.8000 20.2000 45.1000 ;
	    RECT 18.2000 41.1000 18.6000 44.6000 ;
	    RECT 19.8000 41.1000 20.2000 44.8000 ;
	    RECT 20.6000 44.8000 21.7000 45.1000 ;
	    RECT 20.6000 41.1000 21.0000 44.8000 ;
	    RECT 22.2000 41.1000 22.6000 45.1000 ;
	    RECT 23.8000 46.1000 24.2000 49.9000 ;
	    RECT 25.4000 47.8000 25.8000 48.6000 ;
	    RECT 24.6000 46.8000 25.0000 47.6000 ;
	    RECT 25.4000 46.8000 25.8000 47.2000 ;
	    RECT 25.4000 46.1000 25.7000 46.8000 ;
	    RECT 23.8000 45.8000 25.7000 46.1000 ;
	    RECT 23.8000 41.1000 24.2000 45.8000 ;
	    RECT 25.4000 44.1000 25.8000 44.2000 ;
	    RECT 26.2000 44.1000 26.6000 49.9000 ;
	    RECT 27.6000 47.1000 28.0000 49.9000 ;
	    RECT 30.2000 47.9000 30.6000 49.9000 ;
	    RECT 32.3000 48.4000 32.7000 49.9000 ;
	    RECT 32.3000 47.9000 33.0000 48.4000 ;
	    RECT 30.3000 47.8000 30.6000 47.9000 ;
	    RECT 30.3000 47.6000 31.2000 47.8000 ;
	    RECT 30.3000 47.5000 32.4000 47.6000 ;
	    RECT 30.9000 47.3000 32.4000 47.5000 ;
	    RECT 32.0000 47.2000 32.4000 47.3000 ;
	    RECT 27.1000 46.9000 28.0000 47.1000 ;
	    RECT 27.1000 46.8000 27.9000 46.9000 ;
	    RECT 27.1000 45.2000 27.4000 46.8000 ;
	    RECT 30.2000 46.4000 30.6000 47.2000 ;
	    RECT 31.2000 46.9000 31.6000 47.0000 ;
	    RECT 31.1000 46.6000 31.6000 46.9000 ;
	    RECT 31.1000 46.2000 31.4000 46.6000 ;
	    RECT 28.2000 45.8000 29.0000 46.2000 ;
	    RECT 31.0000 45.8000 31.4000 46.2000 ;
	    RECT 27.0000 44.8000 27.4000 45.2000 ;
	    RECT 29.4000 45.1000 29.8000 45.6000 ;
	    RECT 32.0000 45.5000 32.3000 47.2000 ;
	    RECT 32.7000 46.2000 33.0000 47.9000 ;
	    RECT 35.2000 47.1000 35.6000 49.9000 ;
	    RECT 36.6000 47.7000 37.0000 49.9000 ;
	    RECT 38.7000 49.2000 39.3000 49.9000 ;
	    RECT 38.7000 48.9000 39.4000 49.2000 ;
	    RECT 41.0000 48.9000 41.4000 49.9000 ;
	    RECT 43.2000 49.2000 43.6000 49.9000 ;
	    RECT 43.2000 48.9000 44.2000 49.2000 ;
	    RECT 39.0000 48.5000 39.4000 48.9000 ;
	    RECT 41.1000 48.6000 41.4000 48.9000 ;
	    RECT 41.1000 48.3000 42.5000 48.6000 ;
	    RECT 42.1000 48.2000 42.5000 48.3000 ;
	    RECT 43.0000 48.2000 43.4000 48.6000 ;
	    RECT 43.8000 48.5000 44.2000 48.9000 ;
	    RECT 38.1000 47.7000 38.5000 47.8000 ;
	    RECT 36.6000 47.4000 38.5000 47.7000 ;
	    RECT 35.2000 46.9000 36.1000 47.1000 ;
	    RECT 35.3000 46.8000 36.1000 46.9000 ;
	    RECT 32.6000 45.8000 33.0000 46.2000 ;
	    RECT 34.2000 45.8000 35.0000 46.2000 ;
	    RECT 31.1000 45.2000 32.3000 45.5000 ;
	    RECT 30.2000 45.1000 30.6000 45.2000 ;
	    RECT 29.4000 44.8000 30.6000 45.1000 ;
	    RECT 25.4000 43.8000 26.6000 44.1000 ;
	    RECT 26.2000 41.1000 26.6000 43.8000 ;
	    RECT 27.1000 43.5000 27.4000 44.8000 ;
	    RECT 27.8000 43.8000 28.2000 44.6000 ;
	    RECT 27.1000 43.2000 28.9000 43.5000 ;
	    RECT 27.1000 43.1000 27.4000 43.2000 ;
	    RECT 27.0000 41.1000 27.4000 43.1000 ;
	    RECT 28.6000 43.1000 28.9000 43.2000 ;
	    RECT 31.1000 43.1000 31.4000 45.2000 ;
	    RECT 32.7000 45.1000 33.0000 45.8000 ;
	    RECT 28.6000 41.1000 29.0000 43.1000 ;
	    RECT 31.0000 41.1000 31.4000 43.1000 ;
	    RECT 32.6000 44.1000 33.0000 45.1000 ;
	    RECT 33.4000 45.1000 33.8000 45.6000 ;
	    RECT 35.8000 45.2000 36.1000 46.8000 ;
	    RECT 36.6000 45.7000 37.0000 47.4000 ;
	    RECT 40.1000 47.1000 40.5000 47.2000 ;
	    RECT 43.0000 47.1000 43.3000 48.2000 ;
	    RECT 45.4000 47.5000 45.8000 49.9000 ;
	    RECT 47.8000 47.5000 48.2000 49.9000 ;
	    RECT 50.0000 49.2000 50.4000 49.9000 ;
	    RECT 49.4000 48.9000 50.4000 49.2000 ;
	    RECT 52.2000 48.9000 52.6000 49.9000 ;
	    RECT 54.3000 49.2000 54.9000 49.9000 ;
	    RECT 54.2000 48.9000 54.9000 49.2000 ;
	    RECT 49.4000 48.5000 49.8000 48.9000 ;
	    RECT 52.2000 48.6000 52.5000 48.9000 ;
	    RECT 50.2000 48.2000 50.6000 48.6000 ;
	    RECT 51.1000 48.3000 52.5000 48.6000 ;
	    RECT 54.2000 48.5000 54.6000 48.9000 ;
	    RECT 51.1000 48.2000 51.5000 48.3000 ;
	    RECT 44.6000 47.1000 45.4000 47.2000 ;
	    RECT 48.2000 47.1000 49.0000 47.2000 ;
	    RECT 50.3000 47.1000 50.6000 48.2000 ;
	    RECT 55.0000 47.8000 55.4000 48.2000 ;
	    RECT 55.0000 47.7000 55.5000 47.8000 ;
	    RECT 56.6000 47.7000 57.0000 49.9000 ;
	    RECT 55.0000 47.4000 57.0000 47.7000 ;
	    RECT 53.1000 47.1000 53.5000 47.2000 ;
	    RECT 39.9000 46.8000 53.7000 47.1000 ;
	    RECT 39.0000 46.4000 39.4000 46.5000 ;
	    RECT 37.5000 46.1000 39.4000 46.4000 ;
	    RECT 37.5000 46.0000 37.9000 46.1000 ;
	    RECT 38.3000 45.7000 38.7000 45.8000 ;
	    RECT 36.6000 45.4000 38.7000 45.7000 ;
	    RECT 34.2000 45.1000 34.6000 45.2000 ;
	    RECT 33.4000 44.8000 34.6000 45.1000 ;
	    RECT 35.8000 44.8000 36.2000 45.2000 ;
	    RECT 35.0000 44.1000 35.4000 44.6000 ;
	    RECT 32.6000 43.8000 35.4000 44.1000 ;
	    RECT 32.6000 41.1000 33.0000 43.8000 ;
	    RECT 35.8000 43.5000 36.1000 44.8000 ;
	    RECT 34.3000 43.2000 36.1000 43.5000 ;
	    RECT 34.3000 43.1000 34.6000 43.2000 ;
	    RECT 34.2000 41.1000 34.6000 43.1000 ;
	    RECT 35.8000 43.1000 36.1000 43.2000 ;
	    RECT 35.8000 41.1000 36.2000 43.1000 ;
	    RECT 36.6000 41.1000 37.0000 45.4000 ;
	    RECT 39.9000 45.2000 40.2000 46.8000 ;
	    RECT 43.5000 46.7000 43.9000 46.8000 ;
	    RECT 49.7000 46.7000 50.1000 46.8000 ;
	    RECT 43.0000 46.2000 43.4000 46.3000 ;
	    RECT 44.3000 46.2000 44.7000 46.3000 ;
	    RECT 42.2000 45.9000 44.7000 46.2000 ;
	    RECT 48.9000 46.2000 49.3000 46.3000 ;
	    RECT 53.4000 46.2000 53.7000 46.8000 ;
	    RECT 54.2000 46.4000 54.6000 46.5000 ;
	    RECT 48.9000 45.9000 51.4000 46.2000 ;
	    RECT 42.2000 45.8000 42.6000 45.9000 ;
	    RECT 51.0000 45.8000 51.4000 45.9000 ;
	    RECT 53.4000 45.8000 53.8000 46.2000 ;
	    RECT 54.2000 46.1000 56.1000 46.4000 ;
	    RECT 55.7000 46.0000 56.1000 46.1000 ;
	    RECT 43.0000 45.5000 45.8000 45.6000 ;
	    RECT 42.9000 45.4000 45.8000 45.5000 ;
	    RECT 39.0000 44.9000 40.2000 45.2000 ;
	    RECT 40.9000 45.3000 45.8000 45.4000 ;
	    RECT 40.9000 45.1000 43.3000 45.3000 ;
	    RECT 39.0000 44.4000 39.3000 44.9000 ;
	    RECT 38.6000 44.0000 39.3000 44.4000 ;
	    RECT 40.1000 44.5000 40.5000 44.6000 ;
	    RECT 40.9000 44.5000 41.2000 45.1000 ;
	    RECT 40.1000 44.2000 41.2000 44.5000 ;
	    RECT 41.5000 44.5000 44.2000 44.8000 ;
	    RECT 41.5000 44.4000 41.9000 44.5000 ;
	    RECT 43.8000 44.4000 44.2000 44.5000 ;
	    RECT 40.7000 43.7000 41.1000 43.8000 ;
	    RECT 42.1000 43.7000 42.5000 43.8000 ;
	    RECT 39.0000 43.1000 39.4000 43.5000 ;
	    RECT 40.7000 43.4000 42.5000 43.7000 ;
	    RECT 41.1000 43.1000 41.4000 43.4000 ;
	    RECT 43.8000 43.1000 44.2000 43.5000 ;
	    RECT 38.7000 41.1000 39.3000 43.1000 ;
	    RECT 41.0000 41.1000 41.4000 43.1000 ;
	    RECT 43.2000 42.8000 44.2000 43.1000 ;
	    RECT 43.2000 41.1000 43.6000 42.8000 ;
	    RECT 45.4000 41.1000 45.8000 45.3000 ;
	    RECT 47.8000 45.5000 50.6000 45.6000 ;
	    RECT 47.8000 45.4000 50.7000 45.5000 ;
	    RECT 47.8000 45.3000 52.7000 45.4000 ;
	    RECT 47.8000 41.1000 48.2000 45.3000 ;
	    RECT 50.3000 45.1000 52.7000 45.3000 ;
	    RECT 49.4000 44.5000 52.1000 44.8000 ;
	    RECT 49.4000 44.4000 49.8000 44.5000 ;
	    RECT 51.7000 44.4000 52.1000 44.5000 ;
	    RECT 52.4000 44.5000 52.7000 45.1000 ;
	    RECT 53.4000 45.2000 53.7000 45.8000 ;
	    RECT 54.9000 45.7000 55.3000 45.8000 ;
	    RECT 56.6000 45.7000 57.0000 47.4000 ;
	    RECT 57.4000 47.6000 57.8000 49.9000 ;
	    RECT 59.8000 47.6000 60.2000 49.9000 ;
	    RECT 62.2000 47.8000 62.6000 48.6000 ;
	    RECT 57.4000 47.3000 58.5000 47.6000 ;
	    RECT 59.8000 47.3000 60.9000 47.6000 ;
	    RECT 57.4000 45.8000 57.8000 46.6000 ;
	    RECT 58.2000 45.8000 58.5000 47.3000 ;
	    RECT 59.8000 45.8000 60.2000 46.6000 ;
	    RECT 60.6000 45.8000 60.9000 47.3000 ;
	    RECT 54.9000 45.4000 57.0000 45.7000 ;
	    RECT 53.4000 44.9000 54.6000 45.2000 ;
	    RECT 53.1000 44.5000 53.5000 44.6000 ;
	    RECT 52.4000 44.2000 53.5000 44.5000 ;
	    RECT 54.3000 44.4000 54.6000 44.9000 ;
	    RECT 54.3000 44.0000 55.0000 44.4000 ;
	    RECT 51.1000 43.7000 51.5000 43.8000 ;
	    RECT 52.5000 43.7000 52.9000 43.8000 ;
	    RECT 49.4000 43.1000 49.8000 43.5000 ;
	    RECT 51.1000 43.4000 52.9000 43.7000 ;
	    RECT 52.2000 43.1000 52.5000 43.4000 ;
	    RECT 54.2000 43.1000 54.6000 43.5000 ;
	    RECT 49.4000 42.8000 50.4000 43.1000 ;
	    RECT 50.0000 41.1000 50.4000 42.8000 ;
	    RECT 52.2000 41.1000 52.6000 43.1000 ;
	    RECT 54.3000 41.1000 54.9000 43.1000 ;
	    RECT 56.6000 41.1000 57.0000 45.4000 ;
	    RECT 58.2000 45.4000 58.8000 45.8000 ;
	    RECT 60.6000 45.4000 61.2000 45.8000 ;
	    RECT 58.2000 45.1000 58.5000 45.4000 ;
	    RECT 60.6000 45.1000 60.9000 45.4000 ;
	    RECT 57.4000 44.8000 58.5000 45.1000 ;
	    RECT 59.8000 44.8000 60.9000 45.1000 ;
	    RECT 63.0000 45.1000 63.4000 49.9000 ;
	    RECT 64.1000 48.2000 64.5000 49.9000 ;
	    RECT 67.0000 48.9000 67.4000 49.9000 ;
	    RECT 64.1000 47.9000 65.0000 48.2000 ;
	    RECT 63.8000 47.1000 64.2000 47.2000 ;
	    RECT 64.6000 47.1000 65.0000 47.9000 ;
	    RECT 66.2000 47.8000 66.6000 48.6000 ;
	    RECT 67.1000 47.8000 67.4000 48.9000 ;
	    RECT 68.6000 47.9000 69.0000 49.9000 ;
	    RECT 70.7000 48.2000 71.1000 49.9000 ;
	    RECT 63.8000 46.8000 65.0000 47.1000 ;
	    RECT 65.4000 47.1000 65.8000 47.6000 ;
	    RECT 67.1000 47.5000 68.3000 47.8000 ;
	    RECT 67.0000 47.1000 67.5000 47.2000 ;
	    RECT 65.4000 46.8000 67.5000 47.1000 ;
	    RECT 63.8000 45.1000 64.2000 45.2000 ;
	    RECT 63.0000 44.8000 64.2000 45.1000 ;
	    RECT 57.4000 41.1000 57.8000 44.8000 ;
	    RECT 59.8000 41.1000 60.2000 44.8000 ;
	    RECT 63.0000 41.1000 63.4000 44.8000 ;
	    RECT 63.8000 44.4000 64.2000 44.8000 ;
	    RECT 64.6000 41.1000 65.0000 46.8000 ;
	    RECT 67.2000 46.4000 67.6000 46.8000 ;
	    RECT 68.0000 46.0000 68.3000 47.5000 ;
	    RECT 68.7000 46.2000 69.0000 47.9000 ;
	    RECT 70.2000 47.8000 71.3000 48.2000 ;
	    RECT 69.4000 46.8000 69.8000 47.6000 ;
	    RECT 67.9000 45.7000 68.3000 46.0000 ;
	    RECT 68.6000 45.8000 69.0000 46.2000 ;
	    RECT 66.2000 45.6000 68.3000 45.7000 ;
	    RECT 66.2000 45.4000 68.2000 45.6000 ;
	    RECT 66.2000 41.1000 66.6000 45.4000 ;
	    RECT 68.7000 45.2000 69.0000 45.8000 ;
	    RECT 68.6000 45.1000 69.0000 45.2000 ;
	    RECT 68.3000 44.8000 69.0000 45.1000 ;
	    RECT 68.3000 41.1000 68.7000 44.8000 ;
	    RECT 70.2000 41.1000 70.6000 47.8000 ;
	    RECT 71.0000 47.2000 71.3000 47.8000 ;
	    RECT 71.0000 46.8000 71.4000 47.2000 ;
	    RECT 71.0000 45.1000 71.4000 45.2000 ;
	    RECT 71.8000 45.1000 72.2000 49.9000 ;
	    RECT 74.2000 48.9000 74.6000 49.9000 ;
	    RECT 72.6000 47.8000 73.0000 48.6000 ;
	    RECT 73.4000 47.8000 73.8000 48.6000 ;
	    RECT 74.3000 48.1000 74.6000 48.9000 ;
	    RECT 76.6000 48.9000 77.0000 49.9000 ;
	    RECT 79.5000 49.2000 79.9000 49.9000 ;
	    RECT 75.0000 48.1000 75.4000 48.2000 ;
	    RECT 74.2000 47.8000 75.4000 48.1000 ;
	    RECT 74.3000 47.2000 74.6000 47.8000 ;
	    RECT 74.2000 46.8000 74.6000 47.2000 ;
	    RECT 74.3000 45.1000 74.6000 46.8000 ;
	    RECT 76.6000 47.2000 76.9000 48.9000 ;
	    RECT 79.5000 48.8000 80.2000 49.2000 ;
	    RECT 77.4000 47.8000 77.8000 48.6000 ;
	    RECT 79.5000 48.2000 79.9000 48.8000 ;
	    RECT 79.0000 47.9000 79.9000 48.2000 ;
	    RECT 76.6000 47.1000 77.0000 47.2000 ;
	    RECT 78.2000 47.1000 78.6000 47.6000 ;
	    RECT 76.6000 46.8000 78.6000 47.1000 ;
	    RECT 75.0000 45.4000 75.4000 46.2000 ;
	    RECT 75.8000 45.4000 76.2000 46.2000 ;
	    RECT 76.6000 45.1000 76.9000 46.8000 ;
	    RECT 71.0000 44.8000 72.2000 45.1000 ;
	    RECT 71.0000 44.4000 71.4000 44.8000 ;
	    RECT 71.8000 41.1000 72.2000 44.8000 ;
	    RECT 74.2000 44.7000 75.1000 45.1000 ;
	    RECT 74.7000 41.1000 75.1000 44.7000 ;
	    RECT 76.1000 44.7000 77.0000 45.1000 ;
	    RECT 76.1000 41.1000 76.5000 44.7000 ;
	    RECT 79.0000 41.1000 79.4000 47.9000 ;
	    RECT 79.8000 45.1000 80.2000 45.2000 ;
	    RECT 80.6000 45.1000 81.0000 49.9000 ;
	    RECT 83.0000 48.8000 83.4000 49.9000 ;
	    RECT 82.2000 47.8000 82.6000 48.6000 ;
	    RECT 81.4000 46.8000 81.8000 47.6000 ;
	    RECT 83.1000 47.2000 83.4000 48.8000 ;
	    RECT 84.9000 48.2000 85.3000 49.9000 ;
	    RECT 84.9000 47.9000 85.8000 48.2000 ;
	    RECT 87.0000 47.9000 87.4000 49.9000 ;
	    RECT 87.8000 48.0000 88.2000 49.9000 ;
	    RECT 89.4000 48.0000 89.8000 49.9000 ;
	    RECT 87.8000 47.9000 89.8000 48.0000 ;
	    RECT 91.7000 47.9000 92.5000 49.9000 ;
	    RECT 94.2000 47.9000 94.6000 49.9000 ;
	    RECT 95.0000 48.0000 95.4000 49.9000 ;
	    RECT 96.6000 48.0000 97.0000 49.9000 ;
	    RECT 95.0000 47.9000 97.0000 48.0000 ;
	    RECT 83.0000 46.8000 83.4000 47.2000 ;
	    RECT 83.1000 45.1000 83.4000 46.8000 ;
	    RECT 83.8000 45.4000 84.2000 46.2000 ;
	    RECT 79.8000 44.8000 81.0000 45.1000 ;
	    RECT 79.8000 44.4000 80.2000 44.8000 ;
	    RECT 80.6000 41.1000 81.0000 44.8000 ;
	    RECT 83.0000 44.7000 83.9000 45.1000 ;
	    RECT 83.5000 41.1000 83.9000 44.7000 ;
	    RECT 84.6000 44.4000 85.0000 45.2000 ;
	    RECT 85.4000 45.1000 85.8000 47.9000 ;
	    RECT 86.2000 46.8000 86.6000 47.6000 ;
	    RECT 87.1000 47.2000 87.4000 47.9000 ;
	    RECT 87.9000 47.7000 89.7000 47.9000 ;
	    RECT 89.0000 47.2000 89.4000 47.4000 ;
	    RECT 87.0000 46.8000 88.3000 47.2000 ;
	    RECT 89.0000 46.9000 89.8000 47.2000 ;
	    RECT 89.4000 46.8000 89.8000 46.9000 ;
	    RECT 87.0000 45.1000 87.4000 45.2000 ;
	    RECT 88.0000 45.1000 88.3000 46.8000 ;
	    RECT 91.0000 46.4000 91.4000 47.2000 ;
	    RECT 91.9000 46.2000 92.2000 47.9000 ;
	    RECT 94.3000 47.2000 94.6000 47.9000 ;
	    RECT 95.1000 47.7000 96.9000 47.9000 ;
	    RECT 96.2000 47.2000 96.6000 47.4000 ;
	    RECT 94.2000 46.8000 95.5000 47.2000 ;
	    RECT 96.2000 47.1000 97.0000 47.2000 ;
	    RECT 97.4000 47.1000 97.8000 49.9000 ;
	    RECT 101.4000 48.9000 101.8000 49.9000 ;
	    RECT 98.2000 48.1000 98.6000 48.6000 ;
	    RECT 101.4000 48.1000 101.7000 48.9000 ;
	    RECT 98.2000 47.8000 101.7000 48.1000 ;
	    RECT 102.2000 47.8000 102.6000 48.6000 ;
	    RECT 96.2000 46.9000 97.8000 47.1000 ;
	    RECT 90.2000 46.1000 90.6000 46.2000 ;
	    RECT 90.2000 45.8000 91.0000 46.1000 ;
	    RECT 91.8000 45.8000 92.2000 46.2000 ;
	    RECT 90.6000 45.6000 91.0000 45.8000 ;
	    RECT 91.9000 45.7000 92.2000 45.8000 ;
	    RECT 91.9000 45.4000 92.9000 45.7000 ;
	    RECT 93.4000 45.4000 93.8000 46.2000 ;
	    RECT 92.6000 45.1000 92.9000 45.4000 ;
	    RECT 94.2000 45.1000 94.6000 45.2000 ;
	    RECT 95.2000 45.1000 95.5000 46.8000 ;
	    RECT 96.6000 46.8000 97.8000 46.9000 ;
	    RECT 95.8000 45.8000 96.2000 46.6000 ;
	    RECT 96.6000 46.2000 96.9000 46.8000 ;
	    RECT 96.6000 45.8000 97.0000 46.2000 ;
	    RECT 85.4000 44.8000 87.7000 45.1000 ;
	    RECT 88.0000 44.8000 88.5000 45.1000 ;
	    RECT 85.4000 41.1000 85.8000 44.8000 ;
	    RECT 87.4000 44.2000 87.7000 44.8000 ;
	    RECT 88.1000 44.2000 88.5000 44.8000 ;
	    RECT 90.2000 44.8000 92.2000 45.1000 ;
	    RECT 87.4000 43.8000 87.8000 44.2000 ;
	    RECT 88.1000 43.8000 89.0000 44.2000 ;
	    RECT 88.1000 41.1000 88.5000 43.8000 ;
	    RECT 90.2000 41.1000 90.6000 44.8000 ;
	    RECT 91.8000 41.4000 92.2000 44.8000 ;
	    RECT 92.6000 41.7000 93.0000 45.1000 ;
	    RECT 93.4000 41.4000 93.8000 45.1000 ;
	    RECT 94.2000 44.8000 94.9000 45.1000 ;
	    RECT 95.2000 44.8000 95.7000 45.1000 ;
	    RECT 94.6000 44.2000 94.9000 44.8000 ;
	    RECT 95.3000 44.2000 95.7000 44.8000 ;
	    RECT 94.6000 43.8000 95.0000 44.2000 ;
	    RECT 95.3000 43.8000 96.2000 44.2000 ;
	    RECT 91.8000 41.1000 93.8000 41.4000 ;
	    RECT 95.3000 41.1000 95.7000 43.8000 ;
	    RECT 97.4000 41.1000 97.8000 46.8000 ;
	    RECT 101.4000 47.2000 101.7000 47.8000 ;
	    RECT 103.0000 47.7000 103.4000 49.9000 ;
	    RECT 105.1000 49.2000 105.7000 49.9000 ;
	    RECT 105.1000 48.9000 105.8000 49.2000 ;
	    RECT 107.4000 48.9000 107.8000 49.9000 ;
	    RECT 109.6000 49.2000 110.0000 49.9000 ;
	    RECT 109.6000 48.9000 110.6000 49.2000 ;
	    RECT 105.4000 48.5000 105.8000 48.9000 ;
	    RECT 107.5000 48.6000 107.8000 48.9000 ;
	    RECT 107.5000 48.3000 108.9000 48.6000 ;
	    RECT 108.5000 48.2000 108.9000 48.3000 ;
	    RECT 109.4000 48.2000 109.8000 48.6000 ;
	    RECT 110.2000 48.5000 110.6000 48.9000 ;
	    RECT 104.5000 47.7000 104.9000 47.8000 ;
	    RECT 103.0000 47.4000 104.9000 47.7000 ;
	    RECT 101.4000 46.8000 101.8000 47.2000 ;
	    RECT 100.6000 45.4000 101.0000 46.2000 ;
	    RECT 101.4000 45.1000 101.7000 46.8000 ;
	    RECT 103.0000 45.7000 103.4000 47.4000 ;
	    RECT 106.5000 47.1000 106.9000 47.2000 ;
	    RECT 107.8000 47.1000 108.2000 47.2000 ;
	    RECT 109.4000 47.1000 109.7000 48.2000 ;
	    RECT 111.8000 47.5000 112.2000 49.9000 ;
	    RECT 111.0000 47.1000 111.8000 47.2000 ;
	    RECT 106.3000 46.8000 111.8000 47.1000 ;
	    RECT 112.6000 46.8000 113.0000 47.6000 ;
	    RECT 105.4000 46.4000 105.8000 46.5000 ;
	    RECT 103.9000 46.1000 105.8000 46.4000 ;
	    RECT 103.9000 46.0000 104.3000 46.1000 ;
	    RECT 104.7000 45.7000 105.1000 45.8000 ;
	    RECT 103.0000 45.4000 105.1000 45.7000 ;
	    RECT 100.9000 44.7000 101.8000 45.1000 ;
	    RECT 100.9000 41.1000 101.3000 44.7000 ;
	    RECT 103.0000 41.1000 103.4000 45.4000 ;
	    RECT 106.3000 45.2000 106.6000 46.8000 ;
	    RECT 109.9000 46.7000 110.3000 46.8000 ;
	    RECT 110.7000 46.2000 111.1000 46.3000 ;
	    RECT 108.6000 45.9000 111.1000 46.2000 ;
	    RECT 108.6000 45.8000 109.0000 45.9000 ;
	    RECT 109.4000 45.5000 112.2000 45.6000 ;
	    RECT 109.3000 45.4000 112.2000 45.5000 ;
	    RECT 105.4000 44.9000 106.6000 45.2000 ;
	    RECT 107.3000 45.3000 112.2000 45.4000 ;
	    RECT 107.3000 45.1000 109.7000 45.3000 ;
	    RECT 105.4000 44.4000 105.7000 44.9000 ;
	    RECT 105.0000 44.2000 105.7000 44.4000 ;
	    RECT 106.5000 44.5000 106.9000 44.6000 ;
	    RECT 107.3000 44.5000 107.6000 45.1000 ;
	    RECT 106.5000 44.2000 107.6000 44.5000 ;
	    RECT 107.9000 44.5000 110.6000 44.8000 ;
	    RECT 107.9000 44.4000 108.3000 44.5000 ;
	    RECT 110.2000 44.4000 110.6000 44.5000 ;
	    RECT 104.6000 44.0000 105.7000 44.2000 ;
	    RECT 104.6000 43.8000 105.3000 44.0000 ;
	    RECT 107.1000 43.7000 107.5000 43.8000 ;
	    RECT 108.5000 43.7000 108.9000 43.8000 ;
	    RECT 105.4000 43.1000 105.8000 43.5000 ;
	    RECT 107.1000 43.4000 108.9000 43.7000 ;
	    RECT 107.5000 43.1000 107.8000 43.4000 ;
	    RECT 110.2000 43.1000 110.6000 43.5000 ;
	    RECT 105.1000 41.1000 105.7000 43.1000 ;
	    RECT 107.4000 41.1000 107.8000 43.1000 ;
	    RECT 109.6000 42.8000 110.6000 43.1000 ;
	    RECT 109.6000 41.1000 110.0000 42.8000 ;
	    RECT 111.8000 41.1000 112.2000 45.3000 ;
	    RECT 113.4000 41.1000 113.8000 49.9000 ;
	    RECT 114.2000 47.6000 114.6000 49.9000 ;
	    RECT 115.8000 48.2000 116.2000 49.9000 ;
	    RECT 115.8000 47.9000 116.3000 48.2000 ;
	    RECT 114.2000 47.3000 115.5000 47.6000 ;
	    RECT 114.3000 46.2000 114.7000 46.6000 ;
	    RECT 114.2000 45.8000 114.7000 46.2000 ;
	    RECT 115.2000 46.5000 115.5000 47.3000 ;
	    RECT 116.0000 47.2000 116.3000 47.9000 ;
	    RECT 117.4000 47.5000 117.8000 49.9000 ;
	    RECT 119.6000 49.2000 120.0000 49.9000 ;
	    RECT 119.0000 48.9000 120.0000 49.2000 ;
	    RECT 121.8000 48.9000 122.2000 49.9000 ;
	    RECT 123.9000 49.2000 124.5000 49.9000 ;
	    RECT 123.8000 48.9000 124.5000 49.2000 ;
	    RECT 119.0000 48.5000 119.4000 48.9000 ;
	    RECT 121.8000 48.6000 122.1000 48.9000 ;
	    RECT 119.8000 48.2000 120.2000 48.6000 ;
	    RECT 120.7000 48.3000 122.1000 48.6000 ;
	    RECT 123.8000 48.5000 124.2000 48.9000 ;
	    RECT 120.7000 48.2000 121.1000 48.3000 ;
	    RECT 115.8000 46.8000 116.3000 47.2000 ;
	    RECT 117.8000 47.1000 118.6000 47.2000 ;
	    RECT 119.9000 47.1000 120.2000 48.2000 ;
	    RECT 124.7000 47.7000 125.1000 47.8000 ;
	    RECT 126.2000 47.7000 126.6000 49.9000 ;
	    RECT 124.7000 47.4000 126.6000 47.7000 ;
	    RECT 122.7000 47.1000 123.1000 47.2000 ;
	    RECT 117.8000 46.8000 123.3000 47.1000 ;
	    RECT 115.2000 46.1000 115.7000 46.5000 ;
	    RECT 115.2000 45.1000 115.5000 46.1000 ;
	    RECT 116.0000 45.1000 116.3000 46.8000 ;
	    RECT 119.3000 46.7000 119.7000 46.8000 ;
	    RECT 118.5000 46.2000 118.9000 46.3000 ;
	    RECT 118.5000 46.1000 121.0000 46.2000 ;
	    RECT 121.4000 46.1000 121.8000 46.2000 ;
	    RECT 118.5000 45.9000 121.8000 46.1000 ;
	    RECT 120.6000 45.8000 121.8000 45.9000 ;
	    RECT 114.2000 44.8000 115.5000 45.1000 ;
	    RECT 114.2000 41.1000 114.6000 44.8000 ;
	    RECT 115.8000 44.6000 116.3000 45.1000 ;
	    RECT 117.4000 45.5000 120.2000 45.6000 ;
	    RECT 117.4000 45.4000 120.3000 45.5000 ;
	    RECT 117.4000 45.3000 122.3000 45.4000 ;
	    RECT 115.8000 41.1000 116.2000 44.6000 ;
	    RECT 117.4000 41.1000 117.8000 45.3000 ;
	    RECT 119.9000 45.1000 122.3000 45.3000 ;
	    RECT 119.0000 44.5000 121.7000 44.8000 ;
	    RECT 119.0000 44.4000 119.4000 44.5000 ;
	    RECT 121.3000 44.4000 121.7000 44.5000 ;
	    RECT 122.0000 44.5000 122.3000 45.1000 ;
	    RECT 123.0000 45.2000 123.3000 46.8000 ;
	    RECT 123.8000 46.4000 124.2000 46.5000 ;
	    RECT 123.8000 46.1000 125.7000 46.4000 ;
	    RECT 125.3000 46.0000 125.7000 46.1000 ;
	    RECT 124.5000 45.7000 124.9000 45.8000 ;
	    RECT 126.2000 45.7000 126.6000 47.4000 ;
	    RECT 128.6000 47.9000 129.0000 49.9000 ;
	    RECT 131.0000 48.9000 131.4000 49.9000 ;
	    RECT 129.3000 48.2000 129.7000 48.6000 ;
	    RECT 128.6000 47.2000 128.9000 47.9000 ;
	    RECT 129.4000 47.8000 129.8000 48.2000 ;
	    RECT 130.2000 47.8000 130.6000 48.6000 ;
	    RECT 127.8000 46.4000 128.2000 47.2000 ;
	    RECT 128.6000 46.8000 129.0000 47.2000 ;
	    RECT 129.4000 47.1000 129.7000 47.8000 ;
	    RECT 131.1000 47.2000 131.4000 48.9000 ;
	    RECT 132.6000 47.9000 133.0000 49.9000 ;
	    RECT 133.4000 48.0000 133.8000 49.9000 ;
	    RECT 135.0000 48.0000 135.4000 49.9000 ;
	    RECT 133.4000 47.9000 135.4000 48.0000 ;
	    RECT 132.7000 47.2000 133.0000 47.9000 ;
	    RECT 133.5000 47.7000 135.3000 47.9000 ;
	    RECT 135.8000 47.8000 136.2000 48.6000 ;
	    RECT 134.6000 47.2000 135.0000 47.4000 ;
	    RECT 131.0000 47.1000 131.4000 47.2000 ;
	    RECT 129.4000 46.8000 131.4000 47.1000 ;
	    RECT 132.6000 46.8000 133.9000 47.2000 ;
	    RECT 134.6000 46.9000 135.4000 47.2000 ;
	    RECT 135.0000 46.8000 135.4000 46.9000 ;
	    RECT 136.6000 47.1000 137.0000 49.9000 ;
	    RECT 137.4000 48.0000 137.8000 49.9000 ;
	    RECT 139.0000 48.0000 139.4000 49.9000 ;
	    RECT 137.4000 47.9000 139.4000 48.0000 ;
	    RECT 139.8000 47.9000 140.2000 49.9000 ;
	    RECT 137.5000 47.7000 139.3000 47.9000 ;
	    RECT 137.8000 47.2000 138.2000 47.4000 ;
	    RECT 139.8000 47.2000 140.1000 47.9000 ;
	    RECT 140.6000 47.6000 141.0000 49.9000 ;
	    RECT 140.6000 47.3000 141.7000 47.6000 ;
	    RECT 137.4000 47.1000 138.2000 47.2000 ;
	    RECT 136.6000 46.9000 138.2000 47.1000 ;
	    RECT 136.6000 46.8000 137.8000 46.9000 ;
	    RECT 138.9000 46.8000 140.2000 47.2000 ;
	    RECT 127.0000 46.1000 127.4000 46.2000 ;
	    RECT 128.6000 46.1000 128.9000 46.8000 ;
	    RECT 129.4000 46.1000 129.8000 46.2000 ;
	    RECT 127.0000 45.8000 127.8000 46.1000 ;
	    RECT 128.6000 45.8000 129.8000 46.1000 ;
	    RECT 124.5000 45.4000 126.6000 45.7000 ;
	    RECT 127.4000 45.6000 127.8000 45.8000 ;
	    RECT 123.0000 44.9000 124.2000 45.2000 ;
	    RECT 122.7000 44.5000 123.1000 44.6000 ;
	    RECT 122.0000 44.2000 123.1000 44.5000 ;
	    RECT 123.9000 44.4000 124.2000 44.9000 ;
	    RECT 123.9000 44.0000 124.6000 44.4000 ;
	    RECT 120.7000 43.7000 121.1000 43.8000 ;
	    RECT 122.1000 43.7000 122.5000 43.8000 ;
	    RECT 119.0000 43.1000 119.4000 43.5000 ;
	    RECT 120.7000 43.4000 122.5000 43.7000 ;
	    RECT 121.8000 43.1000 122.1000 43.4000 ;
	    RECT 123.8000 43.1000 124.2000 43.5000 ;
	    RECT 119.0000 42.8000 120.0000 43.1000 ;
	    RECT 119.6000 41.1000 120.0000 42.8000 ;
	    RECT 121.8000 41.1000 122.2000 43.1000 ;
	    RECT 123.9000 41.1000 124.5000 43.1000 ;
	    RECT 126.2000 41.1000 126.6000 45.4000 ;
	    RECT 129.4000 45.1000 129.7000 45.8000 ;
	    RECT 131.1000 45.1000 131.4000 46.8000 ;
	    RECT 131.8000 45.4000 132.2000 46.2000 ;
	    RECT 132.6000 45.1000 133.0000 45.2000 ;
	    RECT 133.6000 45.1000 133.9000 46.8000 ;
	    RECT 134.2000 45.8000 134.6000 46.6000 ;
	    RECT 127.0000 44.8000 129.0000 45.1000 ;
	    RECT 127.0000 41.1000 127.4000 44.8000 ;
	    RECT 128.6000 41.1000 129.0000 44.8000 ;
	    RECT 129.4000 41.1000 129.8000 45.1000 ;
	    RECT 131.0000 44.7000 131.9000 45.1000 ;
	    RECT 132.6000 44.8000 133.3000 45.1000 ;
	    RECT 133.6000 44.8000 134.1000 45.1000 ;
	    RECT 131.5000 41.1000 131.9000 44.7000 ;
	    RECT 133.0000 44.2000 133.3000 44.8000 ;
	    RECT 133.0000 43.8000 133.4000 44.2000 ;
	    RECT 133.7000 42.2000 134.1000 44.8000 ;
	    RECT 133.7000 41.8000 134.6000 42.2000 ;
	    RECT 133.7000 41.1000 134.1000 41.8000 ;
	    RECT 136.6000 41.1000 137.0000 46.8000 ;
	    RECT 138.2000 45.8000 138.6000 46.6000 ;
	    RECT 138.9000 45.1000 139.2000 46.8000 ;
	    RECT 140.6000 45.8000 141.0000 46.6000 ;
	    RECT 141.4000 45.8000 141.7000 47.3000 ;
	    RECT 143.0000 46.2000 143.4000 49.9000 ;
	    RECT 144.6000 47.6000 145.0000 49.9000 ;
	    RECT 143.9000 47.3000 145.0000 47.6000 ;
	    RECT 141.4000 45.4000 142.0000 45.8000 ;
	    RECT 139.8000 45.1000 140.2000 45.2000 ;
	    RECT 141.4000 45.1000 141.7000 45.4000 ;
	    RECT 138.7000 44.8000 139.2000 45.1000 ;
	    RECT 139.5000 44.8000 140.2000 45.1000 ;
	    RECT 140.6000 44.8000 141.7000 45.1000 ;
	    RECT 143.0000 45.1000 143.3000 46.2000 ;
	    RECT 143.9000 45.8000 144.2000 47.3000 ;
	    RECT 144.6000 45.8000 145.0000 46.6000 ;
	    RECT 143.6000 45.4000 144.2000 45.8000 ;
	    RECT 143.9000 45.1000 144.2000 45.4000 ;
	    RECT 138.7000 41.1000 139.1000 44.8000 ;
	    RECT 139.5000 44.2000 139.8000 44.8000 ;
	    RECT 139.4000 43.8000 139.8000 44.2000 ;
	    RECT 140.6000 41.1000 141.0000 44.8000 ;
	    RECT 143.0000 41.1000 143.4000 45.1000 ;
	    RECT 143.9000 44.8000 145.0000 45.1000 ;
	    RECT 144.6000 41.1000 145.0000 44.8000 ;
	    RECT 145.4000 41.1000 145.8000 49.9000 ;
	    RECT 2.2000 36.2000 2.6000 39.9000 ;
	    RECT 1.5000 35.9000 2.6000 36.2000 ;
	    RECT 1.5000 35.6000 1.8000 35.9000 ;
	    RECT 1.2000 35.2000 1.8000 35.6000 ;
	    RECT 3.0000 35.6000 3.4000 39.9000 ;
	    RECT 5.1000 37.9000 5.7000 39.9000 ;
	    RECT 7.4000 37.9000 7.8000 39.9000 ;
	    RECT 9.6000 38.2000 10.0000 39.9000 ;
	    RECT 9.6000 37.9000 10.6000 38.2000 ;
	    RECT 5.4000 37.5000 5.8000 37.9000 ;
	    RECT 7.5000 37.6000 7.8000 37.9000 ;
	    RECT 7.1000 37.3000 8.9000 37.6000 ;
	    RECT 10.2000 37.5000 10.6000 37.9000 ;
	    RECT 7.1000 37.2000 7.5000 37.3000 ;
	    RECT 8.5000 37.2000 8.9000 37.3000 ;
	    RECT 5.0000 36.6000 5.7000 37.0000 ;
	    RECT 5.4000 36.1000 5.7000 36.6000 ;
	    RECT 6.5000 36.5000 7.6000 36.8000 ;
	    RECT 6.5000 36.4000 6.9000 36.5000 ;
	    RECT 5.4000 35.8000 6.6000 36.1000 ;
	    RECT 3.0000 35.3000 5.1000 35.6000 ;
	    RECT 1.5000 33.7000 1.8000 35.2000 ;
	    RECT 2.2000 35.1000 2.6000 35.2000 ;
	    RECT 3.0000 35.1000 3.4000 35.3000 ;
	    RECT 4.7000 35.2000 5.1000 35.3000 ;
	    RECT 2.2000 34.8000 3.4000 35.1000 ;
	    RECT 2.2000 34.4000 2.6000 34.8000 ;
	    RECT 1.5000 33.4000 2.6000 33.7000 ;
	    RECT 2.2000 31.1000 2.6000 33.4000 ;
	    RECT 3.0000 33.6000 3.4000 34.8000 ;
	    RECT 3.9000 34.9000 4.3000 35.0000 ;
	    RECT 3.9000 34.6000 5.8000 34.9000 ;
	    RECT 5.4000 34.5000 5.8000 34.6000 ;
	    RECT 6.3000 34.2000 6.6000 35.8000 ;
	    RECT 7.3000 35.9000 7.6000 36.5000 ;
	    RECT 7.9000 36.5000 8.3000 36.6000 ;
	    RECT 10.2000 36.5000 10.6000 36.6000 ;
	    RECT 7.9000 36.2000 10.6000 36.5000 ;
	    RECT 7.3000 35.7000 9.7000 35.9000 ;
	    RECT 11.8000 35.7000 12.2000 39.9000 ;
	    RECT 7.3000 35.6000 12.2000 35.7000 ;
	    RECT 9.3000 35.5000 12.2000 35.6000 ;
	    RECT 9.4000 35.4000 12.2000 35.5000 ;
	    RECT 8.6000 35.1000 9.0000 35.2000 ;
	    RECT 8.6000 34.8000 11.1000 35.1000 ;
	    RECT 9.4000 34.7000 9.8000 34.8000 ;
	    RECT 10.7000 34.7000 11.1000 34.8000 ;
	    RECT 9.9000 34.2000 10.3000 34.3000 ;
	    RECT 6.3000 33.9000 11.8000 34.2000 ;
	    RECT 6.5000 33.8000 6.9000 33.9000 ;
	    RECT 8.6000 33.8000 9.0000 33.9000 ;
	    RECT 3.0000 33.3000 5.0000 33.6000 ;
	    RECT 3.0000 31.1000 3.4000 33.3000 ;
	    RECT 4.5000 33.2000 5.0000 33.3000 ;
	    RECT 4.6000 33.1000 5.0000 33.2000 ;
	    RECT 6.2000 33.1000 6.6000 33.2000 ;
	    RECT 4.6000 32.8000 6.6000 33.1000 ;
	    RECT 9.4000 32.8000 9.7000 33.9000 ;
	    RECT 11.0000 33.8000 11.8000 33.9000 ;
	    RECT 8.5000 32.7000 8.9000 32.8000 ;
	    RECT 5.4000 32.1000 5.8000 32.5000 ;
	    RECT 7.5000 32.4000 8.9000 32.7000 ;
	    RECT 9.4000 32.4000 9.8000 32.8000 ;
	    RECT 7.5000 32.1000 7.8000 32.4000 ;
	    RECT 10.2000 32.1000 10.6000 32.5000 ;
	    RECT 5.1000 31.8000 5.8000 32.1000 ;
	    RECT 5.1000 31.1000 5.7000 31.8000 ;
	    RECT 7.4000 31.1000 7.8000 32.1000 ;
	    RECT 9.6000 31.8000 10.6000 32.1000 ;
	    RECT 9.6000 31.1000 10.0000 31.8000 ;
	    RECT 11.8000 31.1000 12.2000 33.5000 ;
	    RECT 12.6000 32.4000 13.0000 33.2000 ;
	    RECT 13.4000 33.1000 13.8000 39.9000 ;
	    RECT 15.5000 36.3000 15.9000 39.9000 ;
	    RECT 15.0000 35.9000 15.9000 36.3000 ;
	    RECT 15.1000 35.1000 15.4000 35.9000 ;
	    RECT 14.2000 34.8000 15.4000 35.1000 ;
	    RECT 15.8000 34.8000 16.2000 35.6000 ;
	    RECT 14.2000 34.2000 14.5000 34.8000 ;
	    RECT 15.1000 34.2000 15.4000 34.8000 ;
	    RECT 14.2000 33.8000 14.6000 34.2000 ;
	    RECT 15.0000 33.8000 15.4000 34.2000 ;
	    RECT 14.2000 33.1000 14.6000 33.2000 ;
	    RECT 13.4000 32.8000 14.6000 33.1000 ;
	    RECT 13.4000 31.1000 13.8000 32.8000 ;
	    RECT 14.2000 32.4000 14.6000 32.8000 ;
	    RECT 15.1000 32.1000 15.4000 33.8000 ;
	    RECT 16.6000 33.4000 17.0000 34.2000 ;
	    RECT 17.4000 33.1000 17.8000 39.9000 ;
	    RECT 18.2000 35.8000 18.6000 36.6000 ;
	    RECT 19.0000 35.8000 19.4000 36.6000 ;
	    RECT 19.8000 33.1000 20.2000 39.9000 ;
	    RECT 21.4000 37.9000 21.8000 39.9000 ;
	    RECT 21.5000 37.8000 21.8000 37.9000 ;
	    RECT 23.0000 37.9000 23.4000 39.9000 ;
	    RECT 24.7000 39.6000 26.5000 39.9000 ;
	    RECT 24.7000 39.5000 25.0000 39.6000 ;
	    RECT 23.0000 37.8000 23.3000 37.9000 ;
	    RECT 21.5000 37.5000 23.3000 37.8000 ;
	    RECT 21.5000 36.2000 21.8000 37.5000 ;
	    RECT 22.2000 36.4000 22.6000 37.2000 ;
	    RECT 24.6000 36.5000 25.0000 39.5000 ;
	    RECT 26.2000 39.5000 26.5000 39.6000 ;
	    RECT 27.0000 39.6000 29.0000 39.9000 ;
	    RECT 25.4000 36.5000 25.8000 39.3000 ;
	    RECT 26.2000 36.7000 26.6000 39.5000 ;
	    RECT 27.0000 37.0000 27.4000 39.6000 ;
	    RECT 27.8000 36.9000 28.2000 39.3000 ;
	    RECT 28.6000 36.9000 29.0000 39.6000 ;
	    RECT 27.8000 36.7000 28.1000 36.9000 ;
	    RECT 26.2000 36.5000 28.1000 36.7000 ;
	    RECT 25.5000 36.2000 25.8000 36.5000 ;
	    RECT 26.3000 36.4000 28.1000 36.5000 ;
	    RECT 28.7000 36.6000 29.0000 36.9000 ;
	    RECT 30.2000 36.9000 30.6000 39.9000 ;
	    RECT 30.2000 36.6000 30.5000 36.9000 ;
	    RECT 28.7000 36.3000 30.5000 36.6000 ;
	    RECT 32.3000 36.3000 32.7000 39.9000 ;
	    RECT 21.4000 35.8000 21.8000 36.2000 ;
	    RECT 21.5000 34.2000 21.8000 35.8000 ;
	    RECT 23.8000 35.4000 24.2000 36.2000 ;
	    RECT 25.4000 36.1000 25.8000 36.2000 ;
	    RECT 25.4000 35.8000 27.1000 36.1000 ;
	    RECT 31.8000 35.9000 32.7000 36.3000 ;
	    RECT 33.7000 36.3000 34.1000 39.9000 ;
	    RECT 33.7000 35.9000 34.6000 36.3000 ;
	    RECT 22.6000 34.8000 23.4000 35.2000 ;
	    RECT 20.6000 33.4000 21.0000 34.2000 ;
	    RECT 21.5000 34.1000 22.3000 34.2000 ;
	    RECT 21.5000 33.9000 22.4000 34.1000 ;
	    RECT 17.4000 32.8000 18.3000 33.1000 ;
	    RECT 17.9000 32.2000 18.3000 32.8000 ;
	    RECT 19.3000 32.8000 20.2000 33.1000 ;
	    RECT 19.3000 32.2000 19.7000 32.8000 ;
	    RECT 15.0000 31.1000 15.4000 32.1000 ;
	    RECT 17.4000 31.8000 18.3000 32.2000 ;
	    RECT 19.0000 31.8000 19.7000 32.2000 ;
	    RECT 17.9000 31.1000 18.3000 31.8000 ;
	    RECT 19.3000 31.1000 19.7000 31.8000 ;
	    RECT 22.0000 31.1000 22.4000 33.9000 ;
	    RECT 26.8000 32.5000 27.1000 35.8000 ;
	    RECT 27.4000 34.8000 28.2000 35.2000 ;
	    RECT 29.4000 35.1000 29.8000 35.2000 ;
	    RECT 31.0000 35.1000 31.4000 35.2000 ;
	    RECT 29.4000 34.8000 31.4000 35.1000 ;
	    RECT 31.9000 34.2000 32.2000 35.9000 ;
	    RECT 32.6000 34.8000 33.0000 35.6000 ;
	    RECT 33.4000 34.8000 33.8000 35.6000 ;
	    RECT 28.2000 33.8000 29.0000 34.2000 ;
	    RECT 31.8000 34.1000 32.2000 34.2000 ;
	    RECT 29.4000 33.8000 32.2000 34.1000 ;
	    RECT 29.4000 33.2000 29.7000 33.8000 ;
	    RECT 28.9000 32.8000 29.8000 33.2000 ;
	    RECT 26.8000 32.2000 28.8000 32.5000 ;
	    RECT 31.0000 32.4000 31.4000 33.2000 ;
	    RECT 26.8000 32.1000 27.4000 32.2000 ;
	    RECT 27.0000 31.1000 27.4000 32.1000 ;
	    RECT 28.5000 32.1000 28.8000 32.2000 ;
	    RECT 31.9000 32.1000 32.2000 33.8000 ;
	    RECT 34.2000 34.2000 34.5000 35.9000 ;
	    RECT 34.2000 33.8000 34.6000 34.2000 ;
	    RECT 33.4000 33.1000 33.8000 33.2000 ;
	    RECT 34.2000 33.1000 34.5000 33.8000 ;
	    RECT 33.4000 32.8000 34.5000 33.1000 ;
	    RECT 28.5000 31.8000 29.0000 32.1000 ;
	    RECT 28.6000 31.1000 29.0000 31.8000 ;
	    RECT 31.8000 31.1000 32.2000 32.1000 ;
	    RECT 34.2000 32.1000 34.5000 32.8000 ;
	    RECT 35.0000 33.1000 35.4000 33.2000 ;
	    RECT 35.8000 33.1000 36.2000 39.9000 ;
	    RECT 38.7000 36.2000 39.1000 39.9000 ;
	    RECT 39.4000 36.8000 39.8000 37.2000 ;
	    RECT 39.5000 36.2000 39.8000 36.8000 ;
	    RECT 40.9000 36.2000 41.3000 39.9000 ;
	    RECT 38.7000 35.9000 39.2000 36.2000 ;
	    RECT 39.5000 35.9000 40.2000 36.2000 ;
	    RECT 38.8000 35.8000 39.2000 35.9000 ;
	    RECT 39.8000 35.8000 40.2000 35.9000 ;
	    RECT 40.6000 35.9000 41.3000 36.2000 ;
	    RECT 40.6000 35.8000 41.0000 35.9000 ;
	    RECT 37.4000 35.1000 37.8000 35.2000 ;
	    RECT 38.2000 35.1000 38.6000 35.2000 ;
	    RECT 37.4000 34.8000 38.6000 35.1000 ;
	    RECT 38.2000 34.4000 38.6000 34.8000 ;
	    RECT 38.9000 34.2000 39.2000 35.8000 ;
	    RECT 40.6000 35.2000 40.9000 35.8000 ;
	    RECT 43.0000 35.6000 43.4000 39.9000 ;
	    RECT 41.4000 35.4000 43.4000 35.6000 ;
	    RECT 41.3000 35.3000 43.4000 35.4000 ;
	    RECT 40.6000 34.8000 41.0000 35.2000 ;
	    RECT 41.3000 35.0000 41.7000 35.3000 ;
	    RECT 37.4000 34.1000 37.8000 34.2000 ;
	    RECT 37.4000 33.8000 38.2000 34.1000 ;
	    RECT 38.9000 33.8000 40.2000 34.2000 ;
	    RECT 37.8000 33.6000 38.2000 33.8000 ;
	    RECT 37.5000 33.1000 39.3000 33.3000 ;
	    RECT 39.8000 33.1000 40.1000 33.8000 ;
	    RECT 40.6000 33.1000 40.9000 34.8000 ;
	    RECT 41.3000 33.5000 41.6000 35.0000 ;
	    RECT 42.0000 34.2000 42.4000 34.6000 ;
	    RECT 42.1000 33.8000 42.6000 34.2000 ;
	    RECT 41.3000 33.2000 42.5000 33.5000 ;
	    RECT 35.0000 32.8000 36.2000 33.1000 ;
	    RECT 35.0000 32.4000 35.4000 32.8000 ;
	    RECT 34.2000 31.1000 34.6000 32.1000 ;
	    RECT 35.8000 31.1000 36.2000 32.8000 ;
	    RECT 37.4000 33.0000 39.4000 33.1000 ;
	    RECT 37.4000 31.1000 37.8000 33.0000 ;
	    RECT 39.0000 31.1000 39.4000 33.0000 ;
	    RECT 39.8000 31.1000 40.2000 33.1000 ;
	    RECT 40.6000 31.1000 41.0000 33.1000 ;
	    RECT 42.2000 32.1000 42.5000 33.2000 ;
	    RECT 43.0000 32.4000 43.4000 33.2000 ;
	    RECT 44.6000 33.1000 45.0000 39.9000 ;
	    RECT 45.4000 35.8000 45.8000 36.6000 ;
	    RECT 46.2000 35.8000 46.6000 36.2000 ;
	    RECT 47.0000 36.1000 47.4000 39.9000 ;
	    RECT 49.8000 36.8000 50.2000 37.2000 ;
	    RECT 49.8000 36.2000 50.1000 36.8000 ;
	    RECT 50.5000 36.2000 50.9000 39.9000 ;
	    RECT 53.0000 36.8000 53.4000 37.2000 ;
	    RECT 53.0000 36.2000 53.3000 36.8000 ;
	    RECT 53.7000 36.2000 54.1000 39.9000 ;
	    RECT 57.1000 36.3000 57.5000 39.9000 ;
	    RECT 49.4000 36.1000 50.1000 36.2000 ;
	    RECT 47.0000 35.9000 50.1000 36.1000 ;
	    RECT 50.4000 35.9000 50.9000 36.2000 ;
	    RECT 52.6000 35.9000 53.3000 36.2000 ;
	    RECT 53.6000 35.9000 54.1000 36.2000 ;
	    RECT 56.6000 35.9000 57.5000 36.3000 ;
	    RECT 58.6000 36.8000 59.0000 37.2000 ;
	    RECT 58.6000 36.2000 58.9000 36.8000 ;
	    RECT 59.3000 36.2000 59.7000 39.9000 ;
	    RECT 58.2000 35.9000 58.9000 36.2000 ;
	    RECT 59.2000 35.9000 59.7000 36.2000 ;
	    RECT 47.0000 35.8000 49.8000 35.9000 ;
	    RECT 46.2000 35.1000 46.5000 35.8000 ;
	    RECT 47.0000 35.1000 47.4000 35.8000 ;
	    RECT 46.2000 34.8000 47.4000 35.1000 ;
	    RECT 44.6000 32.8000 45.5000 33.1000 ;
	    RECT 45.1000 32.2000 45.5000 32.8000 ;
	    RECT 46.2000 32.4000 46.6000 33.2000 ;
	    RECT 42.2000 31.1000 42.6000 32.1000 ;
	    RECT 44.6000 31.8000 45.5000 32.2000 ;
	    RECT 45.1000 31.1000 45.5000 31.8000 ;
	    RECT 47.0000 31.1000 47.4000 34.8000 ;
	    RECT 50.4000 34.2000 50.7000 35.9000 ;
	    RECT 52.6000 35.8000 53.0000 35.9000 ;
	    RECT 51.0000 35.1000 51.4000 35.2000 ;
	    RECT 51.8000 35.1000 52.2000 35.2000 ;
	    RECT 51.0000 34.8000 52.2000 35.1000 ;
	    RECT 52.6000 35.1000 53.0000 35.2000 ;
	    RECT 53.6000 35.1000 53.9000 35.9000 ;
	    RECT 52.6000 34.8000 53.9000 35.1000 ;
	    RECT 51.0000 34.4000 51.4000 34.8000 ;
	    RECT 53.6000 34.2000 53.9000 34.8000 ;
	    RECT 54.2000 35.1000 54.6000 35.2000 ;
	    RECT 56.7000 35.1000 57.0000 35.9000 ;
	    RECT 58.2000 35.8000 58.6000 35.9000 ;
	    RECT 54.2000 34.8000 57.0000 35.1000 ;
	    RECT 57.4000 34.8000 57.8000 35.6000 ;
	    RECT 54.2000 34.4000 54.6000 34.8000 ;
	    RECT 56.7000 34.2000 57.0000 34.8000 ;
	    RECT 59.2000 34.2000 59.5000 35.9000 ;
	    RECT 59.8000 34.4000 60.2000 35.2000 ;
	    RECT 61.4000 35.1000 61.8000 35.2000 ;
	    RECT 62.2000 35.1000 62.6000 39.9000 ;
	    RECT 61.4000 34.8000 62.6000 35.1000 ;
	    RECT 49.4000 33.8000 50.7000 34.2000 ;
	    RECT 51.8000 34.1000 52.2000 34.2000 ;
	    RECT 51.4000 33.8000 52.2000 34.1000 ;
	    RECT 52.6000 33.8000 53.9000 34.2000 ;
	    RECT 55.0000 34.1000 55.4000 34.2000 ;
	    RECT 54.6000 33.8000 55.4000 34.1000 ;
	    RECT 56.6000 33.8000 57.0000 34.2000 ;
	    RECT 58.2000 33.8000 59.5000 34.2000 ;
	    RECT 60.6000 34.1000 61.0000 34.2000 ;
	    RECT 60.2000 33.8000 61.0000 34.1000 ;
	    RECT 49.5000 33.1000 49.8000 33.8000 ;
	    RECT 51.4000 33.6000 51.8000 33.8000 ;
	    RECT 50.3000 33.1000 52.1000 33.3000 ;
	    RECT 52.7000 33.1000 53.0000 33.8000 ;
	    RECT 54.6000 33.6000 55.0000 33.8000 ;
	    RECT 53.5000 33.1000 55.3000 33.3000 ;
	    RECT 49.4000 31.1000 49.8000 33.1000 ;
	    RECT 50.2000 33.0000 52.2000 33.1000 ;
	    RECT 50.2000 31.1000 50.6000 33.0000 ;
	    RECT 51.8000 31.1000 52.2000 33.0000 ;
	    RECT 52.6000 31.1000 53.0000 33.1000 ;
	    RECT 53.4000 33.0000 55.4000 33.1000 ;
	    RECT 53.4000 31.1000 53.8000 33.0000 ;
	    RECT 55.0000 31.1000 55.4000 33.0000 ;
	    RECT 56.7000 32.1000 57.0000 33.8000 ;
	    RECT 58.3000 33.1000 58.6000 33.8000 ;
	    RECT 60.2000 33.6000 60.6000 33.8000 ;
	    RECT 59.1000 33.1000 60.9000 33.3000 ;
	    RECT 56.6000 31.1000 57.0000 32.1000 ;
	    RECT 58.2000 31.1000 58.6000 33.1000 ;
	    RECT 59.0000 33.0000 61.0000 33.1000 ;
	    RECT 59.0000 31.1000 59.4000 33.0000 ;
	    RECT 60.6000 31.1000 61.0000 33.0000 ;
	    RECT 62.2000 31.1000 62.6000 34.8000 ;
	    RECT 63.0000 33.4000 63.4000 34.2000 ;
	    RECT 63.8000 33.4000 64.2000 34.2000 ;
	    RECT 64.6000 34.1000 65.0000 39.9000 ;
	    RECT 66.2000 36.9000 66.6000 39.9000 ;
	    RECT 66.3000 36.6000 66.6000 36.9000 ;
	    RECT 67.8000 39.6000 69.8000 39.9000 ;
	    RECT 67.8000 36.9000 68.2000 39.6000 ;
	    RECT 68.6000 36.9000 69.0000 39.3000 ;
	    RECT 69.4000 37.0000 69.8000 39.6000 ;
	    RECT 70.3000 39.6000 72.1000 39.9000 ;
	    RECT 70.3000 39.5000 70.6000 39.6000 ;
	    RECT 67.8000 36.6000 68.1000 36.9000 ;
	    RECT 65.4000 35.8000 65.8000 36.6000 ;
	    RECT 66.3000 36.3000 68.1000 36.6000 ;
	    RECT 68.7000 36.7000 69.0000 36.9000 ;
	    RECT 70.2000 36.7000 70.6000 39.5000 ;
	    RECT 71.8000 39.5000 72.1000 39.6000 ;
	    RECT 68.7000 36.5000 70.6000 36.7000 ;
	    RECT 71.0000 36.5000 71.4000 39.3000 ;
	    RECT 71.8000 36.5000 72.2000 39.5000 ;
	    RECT 68.7000 36.4000 70.5000 36.5000 ;
	    RECT 71.0000 36.2000 71.3000 36.5000 ;
	    RECT 71.0000 36.1000 71.4000 36.2000 ;
	    RECT 69.7000 35.8000 71.4000 36.1000 ;
	    RECT 72.6000 35.8000 73.0000 36.6000 ;
	    RECT 68.6000 34.8000 69.4000 35.2000 ;
	    RECT 67.8000 34.1000 68.6000 34.2000 ;
	    RECT 64.6000 33.8000 68.6000 34.1000 ;
	    RECT 64.6000 33.1000 65.0000 33.8000 ;
	    RECT 64.6000 32.8000 65.5000 33.1000 ;
	    RECT 67.0000 32.8000 67.9000 33.2000 ;
	    RECT 65.1000 32.1000 65.5000 32.8000 ;
	    RECT 69.7000 32.5000 70.0000 35.8000 ;
	    RECT 73.4000 33.1000 73.8000 39.9000 ;
	    RECT 75.8000 37.9000 76.2000 39.9000 ;
	    RECT 75.9000 37.8000 76.2000 37.9000 ;
	    RECT 77.4000 37.9000 77.8000 39.9000 ;
	    RECT 77.4000 37.8000 77.7000 37.9000 ;
	    RECT 75.9000 37.5000 77.7000 37.8000 ;
	    RECT 76.6000 36.4000 77.0000 37.2000 ;
	    RECT 77.4000 36.2000 77.7000 37.5000 ;
	    RECT 75.0000 35.4000 75.4000 36.2000 ;
	    RECT 77.4000 35.8000 77.8000 36.2000 ;
	    RECT 75.8000 34.8000 76.6000 35.2000 ;
	    RECT 77.4000 34.2000 77.7000 35.8000 ;
	    RECT 74.2000 33.4000 74.6000 34.2000 ;
	    RECT 76.9000 34.1000 77.7000 34.2000 ;
	    RECT 76.8000 33.9000 77.7000 34.1000 ;
	    RECT 79.0000 34.1000 79.4000 39.9000 ;
	    RECT 79.8000 36.2000 80.2000 39.9000 ;
	    RECT 81.4000 36.2000 81.8000 39.9000 ;
	    RECT 79.8000 35.9000 81.8000 36.2000 ;
	    RECT 82.2000 35.9000 82.6000 39.9000 ;
	    RECT 84.3000 36.3000 84.7000 39.9000 ;
	    RECT 83.8000 35.9000 84.7000 36.3000 ;
	    RECT 80.2000 35.2000 80.6000 35.4000 ;
	    RECT 82.2000 35.2000 82.5000 35.9000 ;
	    RECT 79.8000 34.9000 80.6000 35.2000 ;
	    RECT 81.4000 34.9000 82.6000 35.2000 ;
	    RECT 79.8000 34.8000 80.2000 34.9000 ;
	    RECT 80.6000 34.1000 81.0000 34.6000 ;
	    RECT 68.0000 32.2000 70.0000 32.5000 ;
	    RECT 66.2000 32.1000 66.6000 32.2000 ;
	    RECT 68.0000 32.1000 68.3000 32.2000 ;
	    RECT 65.1000 31.8000 66.6000 32.1000 ;
	    RECT 67.8000 31.8000 68.3000 32.1000 ;
	    RECT 69.4000 32.1000 70.0000 32.2000 ;
	    RECT 71.0000 32.8000 73.8000 33.1000 ;
	    RECT 76.8000 33.1000 77.2000 33.9000 ;
	    RECT 79.0000 33.8000 81.0000 34.1000 ;
	    RECT 78.2000 33.1000 78.6000 33.2000 ;
	    RECT 76.8000 32.8000 78.6000 33.1000 ;
	    RECT 71.0000 32.2000 71.3000 32.8000 ;
	    RECT 65.1000 31.1000 65.5000 31.8000 ;
	    RECT 67.8000 31.1000 68.2000 31.8000 ;
	    RECT 69.4000 31.1000 69.8000 32.1000 ;
	    RECT 71.0000 31.8000 71.4000 32.2000 ;
	    RECT 72.9000 31.1000 73.3000 32.8000 ;
	    RECT 76.8000 31.1000 77.2000 32.8000 ;
	    RECT 78.2000 32.4000 78.6000 32.8000 ;
	    RECT 79.0000 31.1000 79.4000 33.8000 ;
	    RECT 81.4000 33.1000 81.7000 34.9000 ;
	    RECT 82.2000 34.8000 82.6000 34.9000 ;
	    RECT 83.9000 34.2000 84.2000 35.9000 ;
	    RECT 85.4000 35.8000 85.8000 36.6000 ;
	    RECT 84.6000 35.1000 85.0000 35.6000 ;
	    RECT 86.2000 35.1000 86.6000 39.9000 ;
	    RECT 88.1000 36.3000 88.5000 39.9000 ;
	    RECT 90.5000 36.3000 90.9000 39.9000 ;
	    RECT 88.1000 35.9000 89.0000 36.3000 ;
	    RECT 90.5000 35.9000 91.4000 36.3000 ;
	    RECT 84.6000 34.8000 86.6000 35.1000 ;
	    RECT 87.8000 34.8000 88.2000 35.6000 ;
	    RECT 83.8000 34.1000 84.2000 34.2000 ;
	    RECT 82.2000 33.8000 84.2000 34.1000 ;
	    RECT 82.2000 33.2000 82.5000 33.8000 ;
	    RECT 81.4000 31.1000 81.8000 33.1000 ;
	    RECT 82.2000 32.8000 82.6000 33.2000 ;
	    RECT 82.1000 32.4000 82.5000 32.8000 ;
	    RECT 83.0000 32.4000 83.4000 33.2000 ;
	    RECT 83.9000 32.1000 84.2000 33.8000 ;
	    RECT 86.2000 33.1000 86.6000 34.8000 ;
	    RECT 88.6000 34.2000 88.9000 35.9000 ;
	    RECT 90.2000 34.8000 90.6000 35.6000 ;
	    RECT 91.0000 34.2000 91.3000 35.9000 ;
	    RECT 87.0000 34.1000 87.4000 34.2000 ;
	    RECT 88.6000 34.1000 89.0000 34.2000 ;
	    RECT 87.0000 33.8000 89.0000 34.1000 ;
	    RECT 91.0000 34.1000 91.4000 34.2000 ;
	    RECT 91.8000 34.1000 92.2000 34.2000 ;
	    RECT 91.0000 33.8000 92.2000 34.1000 ;
	    RECT 87.0000 33.4000 87.4000 33.8000 ;
	    RECT 83.8000 31.1000 84.2000 32.1000 ;
	    RECT 85.7000 32.8000 86.6000 33.1000 ;
	    RECT 85.7000 31.1000 86.1000 32.8000 ;
	    RECT 88.6000 32.1000 88.9000 33.8000 ;
	    RECT 89.4000 32.4000 89.8000 33.2000 ;
	    RECT 91.0000 32.1000 91.3000 33.8000 ;
	    RECT 91.8000 33.1000 92.2000 33.2000 ;
	    RECT 92.6000 33.1000 93.0000 39.9000 ;
	    RECT 95.0000 36.4000 95.4000 39.9000 ;
	    RECT 94.9000 35.9000 95.4000 36.4000 ;
	    RECT 96.6000 36.2000 97.0000 39.9000 ;
	    RECT 99.8000 36.4000 100.2000 39.9000 ;
	    RECT 95.7000 35.9000 97.0000 36.2000 ;
	    RECT 99.7000 35.9000 100.2000 36.4000 ;
	    RECT 101.4000 36.2000 101.8000 39.9000 ;
	    RECT 100.5000 35.9000 101.8000 36.2000 ;
	    RECT 103.5000 36.2000 103.9000 39.9000 ;
	    RECT 106.2000 37.9000 106.6000 39.9000 ;
	    RECT 104.2000 36.8000 104.6000 37.2000 ;
	    RECT 104.3000 36.2000 104.6000 36.8000 ;
	    RECT 103.5000 35.9000 104.0000 36.2000 ;
	    RECT 104.3000 36.1000 105.0000 36.2000 ;
	    RECT 105.4000 36.1000 105.8000 36.2000 ;
	    RECT 104.3000 35.9000 105.8000 36.1000 ;
	    RECT 94.9000 34.2000 95.2000 35.9000 ;
	    RECT 95.7000 34.9000 96.0000 35.9000 ;
	    RECT 95.5000 34.5000 96.0000 34.9000 ;
	    RECT 94.2000 34.1000 94.6000 34.2000 ;
	    RECT 94.9000 34.1000 95.4000 34.2000 ;
	    RECT 94.2000 33.8000 95.4000 34.1000 ;
	    RECT 91.8000 32.8000 93.0000 33.1000 ;
	    RECT 91.8000 32.4000 92.2000 32.8000 ;
	    RECT 88.6000 31.1000 89.0000 32.1000 ;
	    RECT 91.0000 31.1000 91.4000 32.1000 ;
	    RECT 92.6000 31.1000 93.0000 32.8000 ;
	    RECT 93.4000 32.4000 93.8000 33.2000 ;
	    RECT 94.9000 33.1000 95.2000 33.8000 ;
	    RECT 95.7000 33.7000 96.0000 34.5000 ;
	    RECT 99.7000 34.2000 100.0000 35.9000 ;
	    RECT 100.5000 34.9000 100.8000 35.9000 ;
	    RECT 103.6000 35.8000 104.0000 35.9000 ;
	    RECT 104.6000 35.8000 105.8000 35.9000 ;
	    RECT 106.3000 35.8000 106.6000 37.9000 ;
	    RECT 107.8000 35.9000 108.2000 39.9000 ;
	    RECT 109.9000 36.2000 110.3000 39.9000 ;
	    RECT 110.6000 36.8000 111.0000 37.2000 ;
	    RECT 110.7000 36.2000 111.0000 36.8000 ;
	    RECT 109.9000 35.9000 110.4000 36.2000 ;
	    RECT 110.7000 35.9000 111.4000 36.2000 ;
	    RECT 100.3000 34.5000 100.8000 34.9000 ;
	    RECT 99.0000 34.1000 99.4000 34.2000 ;
	    RECT 99.7000 34.1000 100.2000 34.2000 ;
	    RECT 99.0000 33.8000 100.2000 34.1000 ;
	    RECT 95.7000 33.4000 97.0000 33.7000 ;
	    RECT 94.9000 32.8000 95.4000 33.1000 ;
	    RECT 95.0000 31.1000 95.4000 32.8000 ;
	    RECT 96.6000 31.1000 97.0000 33.4000 ;
	    RECT 99.7000 33.1000 100.0000 33.8000 ;
	    RECT 100.5000 33.7000 100.8000 34.5000 ;
	    RECT 103.0000 34.4000 103.4000 35.2000 ;
	    RECT 103.7000 34.2000 104.0000 35.8000 ;
	    RECT 106.3000 35.5000 107.5000 35.8000 ;
	    RECT 106.2000 34.8000 106.6000 35.2000 ;
	    RECT 102.2000 34.1000 102.6000 34.2000 ;
	    RECT 102.2000 33.8000 103.0000 34.1000 ;
	    RECT 103.7000 33.8000 105.0000 34.2000 ;
	    RECT 105.4000 33.8000 105.8000 34.6000 ;
	    RECT 106.3000 34.4000 106.6000 34.8000 ;
	    RECT 106.3000 34.1000 106.8000 34.4000 ;
	    RECT 106.4000 34.0000 106.8000 34.1000 ;
	    RECT 107.2000 33.8000 107.5000 35.5000 ;
	    RECT 107.9000 35.2000 108.2000 35.9000 ;
	    RECT 110.1000 35.2000 110.4000 35.9000 ;
	    RECT 111.0000 35.8000 111.4000 35.9000 ;
	    RECT 111.8000 35.7000 112.2000 39.9000 ;
	    RECT 114.0000 38.2000 114.4000 39.9000 ;
	    RECT 113.4000 37.9000 114.4000 38.2000 ;
	    RECT 116.2000 37.9000 116.6000 39.9000 ;
	    RECT 118.3000 37.9000 118.9000 39.9000 ;
	    RECT 113.4000 37.5000 113.8000 37.9000 ;
	    RECT 116.2000 37.6000 116.5000 37.9000 ;
	    RECT 115.1000 37.3000 116.9000 37.6000 ;
	    RECT 118.2000 37.5000 118.6000 37.9000 ;
	    RECT 115.1000 37.2000 115.5000 37.3000 ;
	    RECT 116.5000 37.2000 116.9000 37.3000 ;
	    RECT 113.4000 36.5000 113.8000 36.6000 ;
	    RECT 115.7000 36.5000 116.1000 36.6000 ;
	    RECT 113.4000 36.2000 116.1000 36.5000 ;
	    RECT 116.4000 36.5000 117.5000 36.8000 ;
	    RECT 116.4000 35.9000 116.7000 36.5000 ;
	    RECT 117.1000 36.4000 117.5000 36.5000 ;
	    RECT 118.3000 36.6000 119.0000 37.0000 ;
	    RECT 118.3000 36.1000 118.6000 36.6000 ;
	    RECT 114.3000 35.7000 116.7000 35.9000 ;
	    RECT 111.8000 35.6000 116.7000 35.7000 ;
	    RECT 117.4000 35.8000 118.6000 36.1000 ;
	    RECT 111.8000 35.5000 114.7000 35.6000 ;
	    RECT 111.8000 35.4000 114.6000 35.5000 ;
	    RECT 107.8000 35.1000 108.2000 35.2000 ;
	    RECT 107.8000 34.8000 108.9000 35.1000 ;
	    RECT 100.5000 33.4000 101.8000 33.7000 ;
	    RECT 102.6000 33.6000 103.0000 33.8000 ;
	    RECT 99.7000 32.8000 100.2000 33.1000 ;
	    RECT 99.8000 31.1000 100.2000 32.8000 ;
	    RECT 101.4000 31.1000 101.8000 33.4000 ;
	    RECT 102.3000 33.1000 104.1000 33.3000 ;
	    RECT 104.6000 33.1000 104.9000 33.8000 ;
	    RECT 107.2000 33.7000 107.6000 33.8000 ;
	    RECT 106.1000 33.5000 107.6000 33.7000 ;
	    RECT 105.5000 33.4000 107.6000 33.5000 ;
	    RECT 105.5000 33.2000 106.4000 33.4000 ;
	    RECT 105.5000 33.1000 105.8000 33.2000 ;
	    RECT 107.9000 33.1000 108.2000 34.8000 ;
	    RECT 108.6000 34.2000 108.9000 34.8000 ;
	    RECT 109.4000 34.4000 109.8000 35.2000 ;
	    RECT 110.1000 34.8000 110.6000 35.2000 ;
	    RECT 115.0000 35.1000 115.4000 35.2000 ;
	    RECT 112.9000 34.8000 115.4000 35.1000 ;
	    RECT 110.1000 34.2000 110.4000 34.8000 ;
	    RECT 112.9000 34.7000 113.3000 34.8000 ;
	    RECT 114.2000 34.7000 114.6000 34.8000 ;
	    RECT 113.7000 34.2000 114.1000 34.3000 ;
	    RECT 117.4000 34.2000 117.7000 35.8000 ;
	    RECT 120.6000 35.6000 121.0000 39.9000 ;
	    RECT 121.4000 36.2000 121.8000 39.9000 ;
	    RECT 123.0000 36.2000 123.4000 39.9000 ;
	    RECT 121.4000 35.9000 123.4000 36.2000 ;
	    RECT 123.8000 35.9000 124.2000 39.9000 ;
	    RECT 118.9000 35.3000 121.0000 35.6000 ;
	    RECT 118.9000 35.2000 119.3000 35.3000 ;
	    RECT 119.7000 34.9000 120.1000 35.0000 ;
	    RECT 118.2000 34.6000 120.1000 34.9000 ;
	    RECT 118.2000 34.5000 118.6000 34.6000 ;
	    RECT 108.6000 34.1000 109.0000 34.2000 ;
	    RECT 108.6000 33.8000 109.4000 34.1000 ;
	    RECT 110.1000 33.8000 111.4000 34.2000 ;
	    RECT 112.2000 33.9000 117.7000 34.2000 ;
	    RECT 112.2000 33.8000 113.0000 33.9000 ;
	    RECT 109.0000 33.6000 109.4000 33.8000 ;
	    RECT 108.7000 33.1000 110.5000 33.3000 ;
	    RECT 111.0000 33.1000 111.3000 33.8000 ;
	    RECT 102.2000 33.0000 104.2000 33.1000 ;
	    RECT 102.2000 31.1000 102.6000 33.0000 ;
	    RECT 103.8000 31.1000 104.2000 33.0000 ;
	    RECT 104.6000 31.1000 105.0000 33.1000 ;
	    RECT 105.4000 31.1000 105.8000 33.1000 ;
	    RECT 107.5000 32.6000 108.2000 33.1000 ;
	    RECT 108.6000 33.0000 110.6000 33.1000 ;
	    RECT 107.5000 31.1000 107.9000 32.6000 ;
	    RECT 108.6000 31.1000 109.0000 33.0000 ;
	    RECT 110.2000 31.1000 110.6000 33.0000 ;
	    RECT 111.0000 31.1000 111.4000 33.1000 ;
	    RECT 111.8000 31.1000 112.2000 33.5000 ;
	    RECT 114.3000 32.8000 114.6000 33.9000 ;
	    RECT 117.1000 33.8000 117.5000 33.9000 ;
	    RECT 120.6000 33.6000 121.0000 35.3000 ;
	    RECT 121.8000 35.2000 122.2000 35.4000 ;
	    RECT 123.8000 35.2000 124.1000 35.9000 ;
	    RECT 124.6000 35.7000 125.0000 39.9000 ;
	    RECT 126.8000 38.2000 127.2000 39.9000 ;
	    RECT 126.2000 37.9000 127.2000 38.2000 ;
	    RECT 129.0000 37.9000 129.4000 39.9000 ;
	    RECT 131.1000 37.9000 131.7000 39.9000 ;
	    RECT 126.2000 37.5000 126.6000 37.9000 ;
	    RECT 129.0000 37.6000 129.3000 37.9000 ;
	    RECT 127.9000 37.3000 129.7000 37.6000 ;
	    RECT 131.0000 37.5000 131.4000 37.9000 ;
	    RECT 127.9000 37.2000 128.3000 37.3000 ;
	    RECT 129.3000 37.2000 129.7000 37.3000 ;
	    RECT 126.2000 36.5000 126.6000 36.6000 ;
	    RECT 128.5000 36.5000 128.9000 36.6000 ;
	    RECT 126.2000 36.2000 128.9000 36.5000 ;
	    RECT 129.2000 36.5000 130.3000 36.8000 ;
	    RECT 129.2000 35.9000 129.5000 36.5000 ;
	    RECT 129.9000 36.4000 130.3000 36.5000 ;
	    RECT 131.1000 36.6000 131.8000 37.0000 ;
	    RECT 131.1000 36.1000 131.4000 36.6000 ;
	    RECT 127.1000 35.7000 129.5000 35.9000 ;
	    RECT 124.6000 35.6000 129.5000 35.7000 ;
	    RECT 130.2000 35.8000 131.4000 36.1000 ;
	    RECT 124.6000 35.5000 127.5000 35.6000 ;
	    RECT 124.6000 35.4000 127.4000 35.5000 ;
	    RECT 121.4000 34.9000 122.2000 35.2000 ;
	    RECT 123.0000 34.9000 124.2000 35.2000 ;
	    RECT 127.8000 35.1000 128.2000 35.2000 ;
	    RECT 121.4000 34.8000 121.8000 34.9000 ;
	    RECT 122.2000 33.8000 122.6000 34.6000 ;
	    RECT 119.1000 33.3000 121.0000 33.6000 ;
	    RECT 119.1000 33.2000 119.5000 33.3000 ;
	    RECT 113.4000 32.1000 113.8000 32.5000 ;
	    RECT 114.2000 32.4000 114.6000 32.8000 ;
	    RECT 115.1000 32.7000 115.5000 32.8000 ;
	    RECT 115.1000 32.4000 116.5000 32.7000 ;
	    RECT 116.2000 32.1000 116.5000 32.4000 ;
	    RECT 118.2000 32.1000 118.6000 32.5000 ;
	    RECT 113.4000 31.8000 114.4000 32.1000 ;
	    RECT 114.0000 31.1000 114.4000 31.8000 ;
	    RECT 116.2000 31.1000 116.6000 32.1000 ;
	    RECT 118.2000 31.8000 118.9000 32.1000 ;
	    RECT 118.3000 31.1000 118.9000 31.8000 ;
	    RECT 120.6000 31.1000 121.0000 33.3000 ;
	    RECT 123.0000 33.1000 123.3000 34.9000 ;
	    RECT 123.8000 34.8000 124.2000 34.9000 ;
	    RECT 125.7000 34.8000 128.2000 35.1000 ;
	    RECT 125.7000 34.7000 126.1000 34.8000 ;
	    RECT 126.5000 34.2000 126.9000 34.3000 ;
	    RECT 130.2000 34.2000 130.5000 35.8000 ;
	    RECT 133.4000 35.6000 133.8000 39.9000 ;
	    RECT 134.2000 36.2000 134.6000 39.9000 ;
	    RECT 135.8000 36.2000 136.2000 39.9000 ;
	    RECT 134.2000 35.9000 136.2000 36.2000 ;
	    RECT 136.6000 35.9000 137.0000 39.9000 ;
	    RECT 137.7000 36.3000 138.1000 39.9000 ;
	    RECT 137.7000 35.9000 138.6000 36.3000 ;
	    RECT 131.7000 35.3000 133.8000 35.6000 ;
	    RECT 131.7000 35.2000 132.1000 35.3000 ;
	    RECT 132.5000 34.9000 132.9000 35.0000 ;
	    RECT 131.0000 34.6000 132.9000 34.9000 ;
	    RECT 131.0000 34.5000 131.4000 34.6000 ;
	    RECT 125.0000 33.9000 130.5000 34.2000 ;
	    RECT 125.0000 33.8000 125.8000 33.9000 ;
	    RECT 123.0000 31.1000 123.4000 33.1000 ;
	    RECT 123.8000 32.8000 124.2000 33.2000 ;
	    RECT 123.7000 32.4000 124.1000 32.8000 ;
	    RECT 124.6000 31.1000 125.0000 33.5000 ;
	    RECT 127.1000 32.8000 127.4000 33.9000 ;
	    RECT 129.9000 33.8000 130.3000 33.9000 ;
	    RECT 133.4000 33.6000 133.8000 35.3000 ;
	    RECT 134.6000 35.2000 135.0000 35.4000 ;
	    RECT 136.6000 35.2000 136.9000 35.9000 ;
	    RECT 134.2000 34.9000 135.0000 35.2000 ;
	    RECT 135.8000 34.9000 137.0000 35.2000 ;
	    RECT 134.2000 34.8000 134.6000 34.9000 ;
	    RECT 135.0000 33.8000 135.4000 34.6000 ;
	    RECT 131.9000 33.3000 133.8000 33.6000 ;
	    RECT 131.9000 33.2000 132.3000 33.3000 ;
	    RECT 126.2000 32.1000 126.6000 32.5000 ;
	    RECT 127.0000 32.4000 127.4000 32.8000 ;
	    RECT 127.9000 32.7000 128.3000 32.8000 ;
	    RECT 127.9000 32.4000 129.3000 32.7000 ;
	    RECT 129.0000 32.1000 129.3000 32.4000 ;
	    RECT 131.0000 32.1000 131.4000 32.5000 ;
	    RECT 126.2000 31.8000 127.2000 32.1000 ;
	    RECT 126.8000 31.1000 127.2000 31.8000 ;
	    RECT 129.0000 31.1000 129.4000 32.1000 ;
	    RECT 131.0000 31.8000 131.7000 32.1000 ;
	    RECT 131.1000 31.1000 131.7000 31.8000 ;
	    RECT 133.4000 31.1000 133.8000 33.3000 ;
	    RECT 135.8000 33.1000 136.1000 34.9000 ;
	    RECT 136.6000 34.8000 137.0000 34.9000 ;
	    RECT 137.4000 34.8000 137.8000 35.6000 ;
	    RECT 138.2000 34.2000 138.5000 35.9000 ;
	    RECT 138.2000 33.8000 138.6000 34.2000 ;
	    RECT 136.6000 33.1000 137.0000 33.2000 ;
	    RECT 138.2000 33.1000 138.5000 33.8000 ;
	    RECT 135.8000 31.1000 136.2000 33.1000 ;
	    RECT 136.6000 32.8000 138.5000 33.1000 ;
	    RECT 136.5000 32.4000 136.9000 32.8000 ;
	    RECT 138.2000 32.1000 138.5000 32.8000 ;
	    RECT 139.0000 32.4000 139.4000 33.2000 ;
	    RECT 138.2000 31.1000 138.6000 32.1000 ;
	    RECT 139.8000 31.1000 140.2000 39.9000 ;
	    RECT 141.4000 36.2000 141.8000 39.9000 ;
	    RECT 143.8000 36.2000 144.2000 39.9000 ;
	    RECT 141.4000 35.9000 142.5000 36.2000 ;
	    RECT 143.8000 35.9000 144.9000 36.2000 ;
	    RECT 142.2000 35.6000 142.5000 35.9000 ;
	    RECT 144.6000 35.6000 144.9000 35.9000 ;
	    RECT 142.2000 35.2000 142.8000 35.6000 ;
	    RECT 144.6000 35.2000 145.2000 35.6000 ;
	    RECT 141.4000 34.4000 141.8000 35.2000 ;
	    RECT 142.2000 33.7000 142.5000 35.2000 ;
	    RECT 143.8000 34.4000 144.2000 35.2000 ;
	    RECT 144.6000 33.7000 144.9000 35.2000 ;
	    RECT 141.4000 33.4000 142.5000 33.7000 ;
	    RECT 143.8000 33.4000 144.9000 33.7000 ;
	    RECT 140.6000 32.4000 141.0000 33.2000 ;
	    RECT 141.4000 31.1000 141.8000 33.4000 ;
	    RECT 143.8000 31.1000 144.2000 33.4000 ;
	    RECT 0.6000 27.7000 1.0000 29.9000 ;
	    RECT 2.7000 29.2000 3.3000 29.9000 ;
	    RECT 2.7000 28.9000 3.4000 29.2000 ;
	    RECT 5.0000 28.9000 5.4000 29.9000 ;
	    RECT 7.2000 29.2000 7.6000 29.9000 ;
	    RECT 7.2000 28.9000 8.2000 29.2000 ;
	    RECT 3.0000 28.5000 3.4000 28.9000 ;
	    RECT 5.1000 28.6000 5.4000 28.9000 ;
	    RECT 5.1000 28.3000 6.5000 28.6000 ;
	    RECT 6.1000 28.2000 6.5000 28.3000 ;
	    RECT 7.0000 28.2000 7.4000 28.6000 ;
	    RECT 7.8000 28.5000 8.2000 28.9000 ;
	    RECT 2.1000 27.7000 2.5000 27.8000 ;
	    RECT 0.6000 27.4000 2.5000 27.7000 ;
	    RECT 0.6000 25.7000 1.0000 27.4000 ;
	    RECT 4.1000 27.1000 4.5000 27.2000 ;
	    RECT 7.0000 27.1000 7.3000 28.2000 ;
	    RECT 9.4000 27.5000 9.8000 29.9000 ;
	    RECT 10.2000 27.9000 10.6000 29.9000 ;
	    RECT 11.0000 28.0000 11.4000 29.9000 ;
	    RECT 12.6000 28.0000 13.0000 29.9000 ;
	    RECT 11.0000 27.9000 13.0000 28.0000 ;
	    RECT 13.7000 28.2000 14.1000 29.9000 ;
	    RECT 18.2000 28.9000 18.6000 29.9000 ;
	    RECT 19.8000 29.2000 20.2000 29.9000 ;
	    RECT 18.0000 28.8000 18.6000 28.9000 ;
	    RECT 19.7000 28.8000 20.2000 29.2000 ;
	    RECT 18.0000 28.5000 20.0000 28.8000 ;
	    RECT 13.7000 27.9000 14.6000 28.2000 ;
	    RECT 10.3000 27.2000 10.6000 27.9000 ;
	    RECT 11.1000 27.7000 12.9000 27.9000 ;
	    RECT 12.2000 27.2000 12.6000 27.4000 ;
	    RECT 8.6000 27.1000 9.4000 27.2000 ;
	    RECT 3.9000 26.8000 9.4000 27.1000 ;
	    RECT 10.2000 26.8000 11.5000 27.2000 ;
	    RECT 12.2000 27.1000 13.0000 27.2000 ;
	    RECT 14.2000 27.1000 14.6000 27.9000 ;
	    RECT 12.2000 26.9000 14.6000 27.1000 ;
	    RECT 12.6000 26.8000 14.6000 26.9000 ;
	    RECT 15.0000 27.1000 15.4000 27.6000 ;
	    RECT 16.6000 27.1000 17.0000 27.2000 ;
	    RECT 15.0000 26.8000 17.0000 27.1000 ;
	    RECT 3.0000 26.4000 3.4000 26.5000 ;
	    RECT 1.5000 26.1000 3.4000 26.4000 ;
	    RECT 1.5000 26.0000 1.9000 26.1000 ;
	    RECT 2.3000 25.7000 2.7000 25.8000 ;
	    RECT 0.6000 25.4000 2.7000 25.7000 ;
	    RECT 0.6000 21.1000 1.0000 25.4000 ;
	    RECT 3.9000 25.2000 4.2000 26.8000 ;
	    RECT 7.5000 26.7000 7.9000 26.8000 ;
	    RECT 7.0000 26.2000 7.4000 26.3000 ;
	    RECT 8.3000 26.2000 8.7000 26.3000 ;
	    RECT 6.2000 25.9000 8.7000 26.2000 ;
	    RECT 6.2000 25.8000 6.6000 25.9000 ;
	    RECT 7.0000 25.5000 9.8000 25.6000 ;
	    RECT 6.9000 25.4000 9.8000 25.5000 ;
	    RECT 3.0000 24.9000 4.2000 25.2000 ;
	    RECT 4.9000 25.3000 9.8000 25.4000 ;
	    RECT 4.9000 25.1000 7.3000 25.3000 ;
	    RECT 3.0000 24.4000 3.3000 24.9000 ;
	    RECT 2.6000 24.0000 3.3000 24.4000 ;
	    RECT 4.1000 24.5000 4.5000 24.6000 ;
	    RECT 4.9000 24.5000 5.2000 25.1000 ;
	    RECT 4.1000 24.2000 5.2000 24.5000 ;
	    RECT 5.5000 24.5000 8.2000 24.8000 ;
	    RECT 5.5000 24.4000 5.9000 24.5000 ;
	    RECT 7.8000 24.4000 8.2000 24.5000 ;
	    RECT 4.7000 23.7000 5.1000 23.8000 ;
	    RECT 6.1000 23.7000 6.5000 23.8000 ;
	    RECT 3.0000 23.1000 3.4000 23.5000 ;
	    RECT 4.7000 23.4000 6.5000 23.7000 ;
	    RECT 5.1000 23.1000 5.4000 23.4000 ;
	    RECT 7.8000 23.1000 8.2000 23.5000 ;
	    RECT 2.7000 21.1000 3.3000 23.1000 ;
	    RECT 5.0000 21.1000 5.4000 23.1000 ;
	    RECT 7.2000 22.8000 8.2000 23.1000 ;
	    RECT 7.2000 21.1000 7.6000 22.8000 ;
	    RECT 9.4000 21.1000 9.8000 25.3000 ;
	    RECT 10.2000 25.1000 10.6000 25.2000 ;
	    RECT 11.2000 25.1000 11.5000 26.8000 ;
	    RECT 11.8000 25.8000 12.2000 26.6000 ;
	    RECT 10.2000 24.8000 10.9000 25.1000 ;
	    RECT 11.2000 24.8000 11.7000 25.1000 ;
	    RECT 10.6000 24.2000 10.9000 24.8000 ;
	    RECT 10.6000 23.8000 11.0000 24.2000 ;
	    RECT 11.3000 22.2000 11.7000 24.8000 ;
	    RECT 13.4000 24.4000 13.8000 25.2000 ;
	    RECT 11.3000 21.8000 12.2000 22.2000 ;
	    RECT 11.3000 21.1000 11.7000 21.8000 ;
	    RECT 14.2000 21.1000 14.6000 26.8000 ;
	    RECT 18.0000 25.2000 18.3000 28.5000 ;
	    RECT 20.1000 27.8000 21.0000 28.2000 ;
	    RECT 22.2000 28.0000 22.6000 29.9000 ;
	    RECT 23.8000 28.0000 24.2000 29.9000 ;
	    RECT 22.2000 27.9000 24.2000 28.0000 ;
	    RECT 24.6000 27.9000 25.0000 29.9000 ;
	    RECT 26.2000 28.8000 26.6000 29.9000 ;
	    RECT 30.2000 28.9000 30.6000 29.9000 ;
	    RECT 31.8000 29.2000 32.2000 29.9000 ;
	    RECT 30.0000 28.8000 30.6000 28.9000 ;
	    RECT 31.7000 28.9000 32.2000 29.2000 ;
	    RECT 35.0000 28.9000 35.4000 29.9000 ;
	    RECT 31.7000 28.8000 32.0000 28.9000 ;
	    RECT 22.3000 27.7000 24.1000 27.9000 ;
	    RECT 22.6000 27.2000 23.0000 27.4000 ;
	    RECT 24.6000 27.2000 24.9000 27.9000 ;
	    RECT 26.2000 27.2000 26.5000 28.8000 ;
	    RECT 27.0000 27.8000 27.4000 28.6000 ;
	    RECT 30.0000 28.5000 32.0000 28.8000 ;
	    RECT 19.4000 27.1000 20.2000 27.2000 ;
	    RECT 20.6000 27.1000 21.0000 27.2000 ;
	    RECT 19.4000 26.8000 21.0000 27.1000 ;
	    RECT 22.2000 26.9000 23.0000 27.2000 ;
	    RECT 22.2000 26.8000 22.6000 26.9000 ;
	    RECT 23.7000 26.8000 25.0000 27.2000 ;
	    RECT 26.2000 26.8000 26.6000 27.2000 ;
	    RECT 18.6000 26.1000 19.4000 26.2000 ;
	    RECT 19.8000 26.1000 20.2000 26.2000 ;
	    RECT 18.6000 25.8000 20.2000 26.1000 ;
	    RECT 16.6000 24.9000 18.3000 25.2000 ;
	    RECT 23.7000 25.1000 24.0000 26.8000 ;
	    RECT 25.4000 25.4000 25.8000 26.2000 ;
	    RECT 24.6000 25.1000 25.0000 25.2000 ;
	    RECT 26.2000 25.1000 26.5000 26.8000 ;
	    RECT 30.0000 25.2000 30.3000 28.5000 ;
	    RECT 32.1000 28.1000 33.0000 28.2000 ;
	    RECT 35.0000 28.1000 35.3000 28.9000 ;
	    RECT 32.1000 27.8000 35.3000 28.1000 ;
	    RECT 35.8000 27.8000 36.2000 28.6000 ;
	    RECT 38.2000 27.9000 38.6000 29.9000 ;
	    RECT 39.8000 28.0000 40.2000 29.9000 ;
	    RECT 41.4000 29.6000 43.4000 29.9000 ;
	    RECT 41.4000 28.0000 41.8000 29.6000 ;
	    RECT 39.8000 27.9000 41.8000 28.0000 ;
	    RECT 42.2000 27.9000 42.6000 29.3000 ;
	    RECT 43.0000 27.9000 43.4000 29.6000 ;
	    RECT 44.6000 28.9000 45.0000 29.9000 ;
	    RECT 47.8000 29.6000 49.8000 29.9000 ;
	    RECT 35.0000 27.2000 35.3000 27.8000 ;
	    RECT 31.4000 26.8000 32.2000 27.2000 ;
	    RECT 35.0000 26.8000 35.4000 27.2000 ;
	    RECT 36.6000 27.1000 37.0000 27.2000 ;
	    RECT 37.4000 27.1000 37.8000 27.2000 ;
	    RECT 36.6000 26.8000 37.8000 27.1000 ;
	    RECT 30.6000 25.8000 31.4000 26.2000 ;
	    RECT 31.8000 26.1000 32.2000 26.2000 ;
	    RECT 34.2000 26.1000 34.6000 26.2000 ;
	    RECT 31.8000 25.8000 34.6000 26.1000 ;
	    RECT 34.2000 25.4000 34.6000 25.8000 ;
	    RECT 16.6000 24.8000 17.0000 24.9000 ;
	    RECT 16.7000 24.5000 17.0000 24.8000 ;
	    RECT 23.5000 24.8000 24.0000 25.1000 ;
	    RECT 24.3000 24.8000 25.0000 25.1000 ;
	    RECT 17.5000 24.5000 19.3000 24.6000 ;
	    RECT 15.8000 21.5000 16.2000 24.5000 ;
	    RECT 16.6000 21.7000 17.0000 24.5000 ;
	    RECT 17.4000 24.3000 19.3000 24.5000 ;
	    RECT 15.9000 21.4000 16.2000 21.5000 ;
	    RECT 17.4000 21.5000 17.8000 24.3000 ;
	    RECT 19.0000 24.1000 19.3000 24.3000 ;
	    RECT 19.9000 24.4000 21.7000 24.7000 ;
	    RECT 19.9000 24.1000 20.2000 24.4000 ;
	    RECT 17.4000 21.4000 17.7000 21.5000 ;
	    RECT 15.9000 21.1000 17.7000 21.4000 ;
	    RECT 18.2000 21.4000 18.6000 24.0000 ;
	    RECT 19.0000 21.7000 19.4000 24.1000 ;
	    RECT 19.8000 21.4000 20.2000 24.1000 ;
	    RECT 18.2000 21.1000 20.2000 21.4000 ;
	    RECT 21.4000 24.1000 21.7000 24.4000 ;
	    RECT 21.4000 21.1000 21.8000 24.1000 ;
	    RECT 23.5000 21.1000 23.9000 24.8000 ;
	    RECT 24.3000 24.2000 24.6000 24.8000 ;
	    RECT 24.2000 23.8000 24.6000 24.2000 ;
	    RECT 25.7000 24.7000 26.6000 25.1000 ;
	    RECT 28.6000 24.9000 30.3000 25.2000 ;
	    RECT 35.0000 25.1000 35.3000 26.8000 ;
	    RECT 37.4000 26.4000 37.8000 26.8000 ;
	    RECT 38.2000 27.1000 38.5000 27.9000 ;
	    RECT 39.9000 27.7000 41.7000 27.9000 ;
	    RECT 40.2000 27.2000 40.6000 27.4000 ;
	    RECT 42.3000 27.2000 42.6000 27.9000 ;
	    RECT 44.6000 27.2000 44.9000 28.9000 ;
	    RECT 45.4000 27.8000 45.8000 28.6000 ;
	    RECT 47.8000 27.9000 48.2000 29.6000 ;
	    RECT 48.6000 27.9000 49.0000 29.3000 ;
	    RECT 49.4000 28.0000 49.8000 29.6000 ;
	    RECT 51.0000 28.0000 51.4000 29.9000 ;
	    RECT 49.4000 27.9000 51.4000 28.0000 ;
	    RECT 52.6000 28.9000 53.0000 29.9000 ;
	    RECT 48.6000 27.2000 48.9000 27.9000 ;
	    RECT 49.5000 27.7000 51.3000 27.9000 ;
	    RECT 50.6000 27.2000 51.0000 27.4000 ;
	    RECT 52.6000 27.2000 52.9000 28.9000 ;
	    RECT 53.4000 27.8000 53.8000 28.6000 ;
	    RECT 39.0000 27.1000 39.4000 27.2000 ;
	    RECT 38.2000 26.8000 39.4000 27.1000 ;
	    RECT 39.8000 26.9000 40.6000 27.2000 ;
	    RECT 41.4000 26.9000 42.6000 27.2000 ;
	    RECT 43.0000 27.1000 43.4000 27.2000 ;
	    RECT 43.8000 27.1000 44.2000 27.2000 ;
	    RECT 39.8000 26.8000 40.2000 26.9000 ;
	    RECT 41.4000 26.8000 41.8000 26.9000 ;
	    RECT 43.0000 26.8000 44.2000 27.1000 ;
	    RECT 44.6000 26.8000 45.0000 27.2000 ;
	    RECT 38.2000 26.1000 38.5000 26.8000 ;
	    RECT 39.0000 26.1000 39.4000 26.2000 ;
	    RECT 38.2000 25.8000 39.4000 26.1000 ;
	    RECT 40.6000 25.8000 41.0000 26.6000 ;
	    RECT 39.0000 25.1000 39.3000 25.8000 ;
	    RECT 41.4000 25.1000 41.7000 26.8000 ;
	    RECT 42.2000 25.8000 42.6000 26.6000 ;
	    RECT 43.0000 26.1000 43.4000 26.8000 ;
	    RECT 43.8000 26.1000 44.2000 26.2000 ;
	    RECT 43.0000 25.8000 44.2000 26.1000 ;
	    RECT 43.8000 25.4000 44.2000 25.8000 ;
	    RECT 44.6000 26.1000 44.9000 26.8000 ;
	    RECT 47.8000 26.4000 48.2000 27.2000 ;
	    RECT 48.6000 26.9000 49.8000 27.2000 ;
	    RECT 50.6000 27.1000 51.4000 27.2000 ;
	    RECT 51.8000 27.1000 52.2000 27.2000 ;
	    RECT 50.6000 26.9000 52.2000 27.1000 ;
	    RECT 49.4000 26.8000 49.8000 26.9000 ;
	    RECT 51.0000 26.8000 52.2000 26.9000 ;
	    RECT 52.6000 26.8000 53.0000 27.2000 ;
	    RECT 53.4000 27.1000 53.8000 27.2000 ;
	    RECT 54.8000 27.1000 55.2000 29.9000 ;
	    RECT 57.4000 27.9000 57.8000 29.9000 ;
	    RECT 58.2000 28.0000 58.6000 29.9000 ;
	    RECT 59.8000 28.0000 60.2000 29.9000 ;
	    RECT 58.2000 27.9000 60.2000 28.0000 ;
	    RECT 61.4000 28.9000 61.8000 29.9000 ;
	    RECT 57.5000 27.2000 57.8000 27.9000 ;
	    RECT 58.3000 27.7000 60.1000 27.9000 ;
	    RECT 59.4000 27.2000 59.8000 27.4000 ;
	    RECT 61.4000 27.2000 61.7000 28.9000 ;
	    RECT 53.4000 26.9000 55.2000 27.1000 ;
	    RECT 53.4000 26.8000 55.1000 26.9000 ;
	    RECT 57.4000 26.8000 58.7000 27.2000 ;
	    RECT 59.4000 26.9000 60.2000 27.2000 ;
	    RECT 59.8000 26.8000 60.2000 26.9000 ;
	    RECT 61.4000 26.8000 61.8000 27.2000 ;
	    RECT 63.6000 27.1000 64.0000 29.9000 ;
	    RECT 67.8000 29.2000 68.2000 29.9000 ;
	    RECT 67.8000 28.9000 68.3000 29.2000 ;
	    RECT 68.0000 28.8000 68.3000 28.9000 ;
	    RECT 69.4000 28.9000 69.8000 29.9000 ;
	    RECT 69.4000 28.8000 70.0000 28.9000 ;
	    RECT 68.0000 28.5000 70.0000 28.8000 ;
	    RECT 66.2000 28.1000 66.6000 28.2000 ;
	    RECT 67.0000 28.1000 67.9000 28.2000 ;
	    RECT 66.2000 27.8000 67.9000 28.1000 ;
	    RECT 63.1000 26.9000 64.0000 27.1000 ;
	    RECT 63.1000 26.8000 63.9000 26.9000 ;
	    RECT 67.8000 26.8000 68.6000 27.2000 ;
	    RECT 45.4000 26.1000 45.8000 26.2000 ;
	    RECT 44.6000 25.8000 45.8000 26.1000 ;
	    RECT 48.6000 25.8000 49.0000 26.6000 ;
	    RECT 44.6000 25.1000 44.9000 25.8000 ;
	    RECT 49.5000 25.2000 49.8000 26.8000 ;
	    RECT 50.2000 26.1000 50.6000 26.6000 ;
	    RECT 51.0000 26.1000 51.4000 26.2000 ;
	    RECT 50.2000 25.8000 51.4000 26.1000 ;
	    RECT 51.8000 25.4000 52.2000 26.2000 ;
	    RECT 52.6000 26.1000 52.9000 26.8000 ;
	    RECT 53.4000 26.1000 53.8000 26.2000 ;
	    RECT 52.6000 25.8000 53.8000 26.1000 ;
	    RECT 49.5000 25.1000 50.6000 25.2000 ;
	    RECT 52.6000 25.1000 52.9000 25.8000 ;
	    RECT 54.3000 25.2000 54.6000 26.8000 ;
	    RECT 55.4000 25.8000 56.2000 26.2000 ;
	    RECT 57.4000 26.1000 57.8000 26.2000 ;
	    RECT 58.4000 26.1000 58.7000 26.8000 ;
	    RECT 57.4000 25.8000 58.7000 26.1000 ;
	    RECT 59.0000 25.8000 59.4000 26.6000 ;
	    RECT 28.6000 24.8000 29.0000 24.9000 ;
	    RECT 25.7000 21.1000 26.1000 24.7000 ;
	    RECT 28.7000 24.5000 29.0000 24.8000 ;
	    RECT 34.5000 24.7000 35.4000 25.1000 ;
	    RECT 36.6000 24.8000 38.6000 25.1000 ;
	    RECT 29.5000 24.5000 31.3000 24.6000 ;
	    RECT 27.8000 21.5000 28.2000 24.5000 ;
	    RECT 28.6000 21.7000 29.0000 24.5000 ;
	    RECT 29.4000 24.3000 31.3000 24.5000 ;
	    RECT 27.9000 21.4000 28.2000 21.5000 ;
	    RECT 29.4000 21.5000 29.8000 24.3000 ;
	    RECT 31.0000 24.1000 31.3000 24.3000 ;
	    RECT 31.9000 24.4000 33.7000 24.7000 ;
	    RECT 31.9000 24.1000 32.2000 24.4000 ;
	    RECT 29.4000 21.4000 29.7000 21.5000 ;
	    RECT 27.9000 21.1000 29.7000 21.4000 ;
	    RECT 30.2000 21.4000 30.6000 24.0000 ;
	    RECT 31.0000 21.7000 31.4000 24.1000 ;
	    RECT 31.8000 21.4000 32.2000 24.1000 ;
	    RECT 30.2000 21.1000 32.2000 21.4000 ;
	    RECT 33.4000 24.1000 33.7000 24.4000 ;
	    RECT 33.4000 21.1000 33.8000 24.1000 ;
	    RECT 34.5000 21.1000 34.9000 24.7000 ;
	    RECT 36.6000 21.1000 37.0000 24.8000 ;
	    RECT 38.2000 21.1000 38.6000 24.8000 ;
	    RECT 39.0000 21.1000 39.4000 25.1000 ;
	    RECT 41.1000 21.1000 42.1000 25.1000 ;
	    RECT 44.1000 24.7000 45.0000 25.1000 ;
	    RECT 49.1000 24.8000 50.6000 25.1000 ;
	    RECT 44.1000 21.1000 44.5000 24.7000 ;
	    RECT 49.1000 21.1000 50.1000 24.8000 ;
	    RECT 52.1000 24.7000 53.0000 25.1000 ;
	    RECT 54.2000 24.8000 54.6000 25.2000 ;
	    RECT 56.6000 24.8000 57.0000 25.6000 ;
	    RECT 58.4000 25.1000 58.7000 25.8000 ;
	    RECT 60.6000 25.4000 61.0000 26.2000 ;
	    RECT 61.4000 25.2000 61.7000 26.8000 ;
	    RECT 63.1000 25.2000 63.4000 26.8000 ;
	    RECT 64.2000 25.8000 65.0000 26.2000 ;
	    RECT 68.6000 25.8000 69.4000 26.2000 ;
	    RECT 61.4000 25.1000 61.8000 25.2000 ;
	    RECT 58.4000 24.8000 58.9000 25.1000 ;
	    RECT 52.1000 21.1000 52.5000 24.7000 ;
	    RECT 54.3000 23.5000 54.6000 24.8000 ;
	    RECT 55.0000 23.8000 55.4000 24.6000 ;
	    RECT 54.3000 23.2000 56.1000 23.5000 ;
	    RECT 54.3000 23.1000 54.6000 23.2000 ;
	    RECT 54.2000 21.1000 54.6000 23.1000 ;
	    RECT 55.8000 23.1000 56.1000 23.2000 ;
	    RECT 55.8000 21.1000 56.2000 23.1000 ;
	    RECT 58.5000 21.1000 58.9000 24.8000 ;
	    RECT 60.9000 24.7000 61.8000 25.1000 ;
	    RECT 63.0000 24.8000 63.4000 25.2000 ;
	    RECT 65.4000 24.8000 65.8000 25.6000 ;
	    RECT 69.7000 25.2000 70.0000 28.5000 ;
	    RECT 71.8000 27.1000 72.2000 27.2000 ;
	    RECT 72.6000 27.1000 73.0000 27.6000 ;
	    RECT 71.8000 26.8000 73.0000 27.1000 ;
	    RECT 72.6000 26.1000 73.0000 26.2000 ;
	    RECT 73.4000 26.1000 73.8000 29.9000 ;
	    RECT 74.2000 27.9000 74.6000 29.9000 ;
	    RECT 75.0000 28.0000 75.4000 29.9000 ;
	    RECT 76.6000 28.0000 77.0000 29.9000 ;
	    RECT 75.0000 27.9000 77.0000 28.0000 ;
	    RECT 78.2000 28.9000 78.6000 29.9000 ;
	    RECT 74.3000 27.2000 74.6000 27.9000 ;
	    RECT 75.1000 27.7000 76.9000 27.9000 ;
	    RECT 76.2000 27.2000 76.6000 27.4000 ;
	    RECT 78.2000 27.2000 78.5000 28.9000 ;
	    RECT 79.0000 27.8000 79.4000 28.6000 ;
	    RECT 79.8000 27.9000 80.2000 29.9000 ;
	    RECT 81.9000 28.4000 82.3000 29.9000 ;
	    RECT 81.9000 27.9000 82.6000 28.4000 ;
	    RECT 79.9000 27.8000 80.2000 27.9000 ;
	    RECT 79.9000 27.6000 80.8000 27.8000 ;
	    RECT 79.9000 27.5000 82.0000 27.6000 ;
	    RECT 80.5000 27.3000 82.0000 27.5000 ;
	    RECT 81.6000 27.2000 82.0000 27.3000 ;
	    RECT 74.2000 26.8000 75.5000 27.2000 ;
	    RECT 76.2000 26.9000 77.0000 27.2000 ;
	    RECT 76.6000 26.8000 77.0000 26.9000 ;
	    RECT 78.2000 26.8000 78.6000 27.2000 ;
	    RECT 72.6000 25.8000 73.8000 26.1000 ;
	    RECT 69.7000 24.9000 71.4000 25.2000 ;
	    RECT 71.0000 24.8000 71.4000 24.9000 ;
	    RECT 73.4000 25.1000 73.8000 25.8000 ;
	    RECT 75.2000 25.2000 75.5000 26.8000 ;
	    RECT 75.8000 25.8000 76.2000 26.6000 ;
	    RECT 76.6000 26.1000 77.0000 26.2000 ;
	    RECT 77.4000 26.1000 77.8000 26.2000 ;
	    RECT 76.6000 25.8000 77.8000 26.1000 ;
	    RECT 77.4000 25.4000 77.8000 25.8000 ;
	    RECT 74.2000 25.1000 74.6000 25.2000 ;
	    RECT 73.4000 24.8000 74.9000 25.1000 ;
	    RECT 75.2000 24.8000 76.2000 25.2000 ;
	    RECT 78.2000 25.1000 78.5000 26.8000 ;
	    RECT 79.8000 26.4000 80.2000 27.2000 ;
	    RECT 80.8000 26.9000 81.2000 27.0000 ;
	    RECT 80.7000 26.6000 81.2000 26.9000 ;
	    RECT 80.7000 26.2000 81.0000 26.6000 ;
	    RECT 80.6000 25.8000 81.0000 26.2000 ;
	    RECT 81.6000 25.5000 81.9000 27.2000 ;
	    RECT 82.3000 26.2000 82.6000 27.9000 ;
	    RECT 82.2000 25.8000 82.6000 26.2000 ;
	    RECT 80.7000 25.2000 81.9000 25.5000 ;
	    RECT 82.3000 25.2000 82.6000 25.8000 ;
	    RECT 60.9000 21.1000 61.3000 24.7000 ;
	    RECT 63.1000 23.5000 63.4000 24.8000 ;
	    RECT 63.8000 23.8000 64.2000 24.6000 ;
	    RECT 66.3000 24.4000 68.1000 24.7000 ;
	    RECT 66.3000 24.1000 66.6000 24.4000 ;
	    RECT 63.1000 23.2000 64.9000 23.5000 ;
	    RECT 63.1000 23.1000 63.4000 23.2000 ;
	    RECT 63.0000 21.1000 63.4000 23.1000 ;
	    RECT 64.6000 23.1000 64.9000 23.2000 ;
	    RECT 64.6000 21.1000 65.0000 23.1000 ;
	    RECT 66.2000 21.1000 66.6000 24.1000 ;
	    RECT 67.8000 24.1000 68.1000 24.4000 ;
	    RECT 68.7000 24.5000 70.5000 24.6000 ;
	    RECT 71.0000 24.5000 71.3000 24.8000 ;
	    RECT 68.7000 24.3000 70.6000 24.5000 ;
	    RECT 68.7000 24.1000 69.0000 24.3000 ;
	    RECT 67.8000 21.4000 68.2000 24.1000 ;
	    RECT 68.6000 21.7000 69.0000 24.1000 ;
	    RECT 69.4000 21.4000 69.8000 24.0000 ;
	    RECT 70.2000 21.5000 70.6000 24.3000 ;
	    RECT 71.0000 21.7000 71.4000 24.5000 ;
	    RECT 67.8000 21.1000 69.8000 21.4000 ;
	    RECT 70.3000 21.4000 70.6000 21.5000 ;
	    RECT 71.8000 21.5000 72.2000 24.5000 ;
	    RECT 71.8000 21.4000 72.1000 21.5000 ;
	    RECT 70.3000 21.1000 72.1000 21.4000 ;
	    RECT 73.4000 21.1000 73.8000 24.8000 ;
	    RECT 74.6000 24.2000 74.9000 24.8000 ;
	    RECT 74.6000 23.8000 75.0000 24.2000 ;
	    RECT 75.3000 21.1000 75.7000 24.8000 ;
	    RECT 77.7000 24.7000 78.6000 25.1000 ;
	    RECT 77.7000 22.2000 78.1000 24.7000 ;
	    RECT 80.7000 23.1000 81.0000 25.2000 ;
	    RECT 77.4000 21.8000 78.1000 22.2000 ;
	    RECT 77.7000 21.1000 78.1000 21.8000 ;
	    RECT 80.6000 21.1000 81.0000 23.1000 ;
	    RECT 82.2000 21.1000 82.6000 25.2000 ;
	    RECT 83.0000 21.1000 83.4000 29.9000 ;
	    RECT 83.8000 28.1000 84.2000 28.6000 ;
	    RECT 84.9000 28.2000 85.3000 29.9000 ;
	    RECT 84.9000 28.1000 85.8000 28.2000 ;
	    RECT 83.8000 27.8000 85.8000 28.1000 ;
	    RECT 84.6000 24.4000 85.0000 25.2000 ;
	    RECT 85.4000 21.1000 85.8000 27.8000 ;
	    RECT 86.2000 26.8000 86.6000 27.6000 ;
	    RECT 87.0000 26.8000 87.4000 27.6000 ;
	    RECT 87.8000 21.1000 88.2000 29.9000 ;
	    RECT 88.6000 27.5000 89.0000 29.9000 ;
	    RECT 90.8000 29.2000 91.2000 29.9000 ;
	    RECT 90.2000 28.9000 91.2000 29.2000 ;
	    RECT 93.0000 28.9000 93.4000 29.9000 ;
	    RECT 95.1000 29.2000 95.7000 29.9000 ;
	    RECT 95.0000 28.9000 95.7000 29.2000 ;
	    RECT 97.4000 29.1000 97.8000 29.9000 ;
	    RECT 98.2000 29.1000 98.6000 29.2000 ;
	    RECT 90.2000 28.5000 90.6000 28.9000 ;
	    RECT 93.0000 28.6000 93.3000 28.9000 ;
	    RECT 91.0000 28.2000 91.4000 28.6000 ;
	    RECT 91.9000 28.3000 93.3000 28.6000 ;
	    RECT 95.0000 28.5000 95.4000 28.9000 ;
	    RECT 97.4000 28.8000 98.6000 29.1000 ;
	    RECT 91.9000 28.2000 92.3000 28.3000 ;
	    RECT 89.0000 27.1000 89.8000 27.2000 ;
	    RECT 91.1000 27.1000 91.4000 28.2000 ;
	    RECT 95.9000 27.7000 96.3000 27.8000 ;
	    RECT 97.4000 27.7000 97.8000 28.8000 ;
	    RECT 95.9000 27.4000 97.8000 27.7000 ;
	    RECT 93.9000 27.1000 94.3000 27.2000 ;
	    RECT 89.0000 26.8000 94.5000 27.1000 ;
	    RECT 90.5000 26.7000 90.9000 26.8000 ;
	    RECT 89.7000 26.2000 90.1000 26.3000 ;
	    RECT 94.2000 26.2000 94.5000 26.8000 ;
	    RECT 95.0000 26.4000 95.4000 26.5000 ;
	    RECT 89.7000 25.9000 92.2000 26.2000 ;
	    RECT 91.8000 25.8000 92.2000 25.9000 ;
	    RECT 94.2000 25.8000 94.6000 26.2000 ;
	    RECT 95.0000 26.1000 96.9000 26.4000 ;
	    RECT 96.5000 26.0000 96.9000 26.1000 ;
	    RECT 88.6000 25.5000 91.4000 25.6000 ;
	    RECT 88.6000 25.4000 91.5000 25.5000 ;
	    RECT 88.6000 25.3000 93.5000 25.4000 ;
	    RECT 88.6000 21.1000 89.0000 25.3000 ;
	    RECT 91.1000 25.1000 93.5000 25.3000 ;
	    RECT 90.2000 24.5000 92.9000 24.8000 ;
	    RECT 90.2000 24.4000 90.6000 24.5000 ;
	    RECT 92.5000 24.4000 92.9000 24.5000 ;
	    RECT 93.2000 24.5000 93.5000 25.1000 ;
	    RECT 94.2000 25.2000 94.5000 25.8000 ;
	    RECT 95.7000 25.7000 96.1000 25.8000 ;
	    RECT 97.4000 25.7000 97.8000 27.4000 ;
	    RECT 99.8000 27.6000 100.2000 29.9000 ;
	    RECT 102.2000 27.6000 102.6000 29.9000 ;
	    RECT 104.6000 27.7000 105.0000 29.9000 ;
	    RECT 106.7000 29.2000 107.3000 29.9000 ;
	    RECT 106.7000 28.9000 107.4000 29.2000 ;
	    RECT 109.0000 28.9000 109.4000 29.9000 ;
	    RECT 111.2000 29.2000 111.6000 29.9000 ;
	    RECT 111.2000 28.9000 112.2000 29.2000 ;
	    RECT 107.0000 28.5000 107.4000 28.9000 ;
	    RECT 109.1000 28.6000 109.4000 28.9000 ;
	    RECT 109.1000 28.3000 110.5000 28.6000 ;
	    RECT 110.1000 28.2000 110.5000 28.3000 ;
	    RECT 111.0000 28.2000 111.4000 28.6000 ;
	    RECT 111.8000 28.5000 112.2000 28.9000 ;
	    RECT 106.1000 27.7000 106.5000 27.8000 ;
	    RECT 99.8000 27.3000 100.9000 27.6000 ;
	    RECT 102.2000 27.3000 103.3000 27.6000 ;
	    RECT 98.2000 26.1000 98.6000 26.2000 ;
	    RECT 99.8000 26.1000 100.2000 26.6000 ;
	    RECT 98.2000 25.8000 100.2000 26.1000 ;
	    RECT 100.6000 25.8000 100.9000 27.3000 ;
	    RECT 102.2000 25.8000 102.6000 26.6000 ;
	    RECT 103.0000 25.8000 103.3000 27.3000 ;
	    RECT 104.6000 27.4000 106.5000 27.7000 ;
	    RECT 95.7000 25.4000 97.8000 25.7000 ;
	    RECT 94.2000 24.9000 95.4000 25.2000 ;
	    RECT 93.9000 24.5000 94.3000 24.6000 ;
	    RECT 93.2000 24.2000 94.3000 24.5000 ;
	    RECT 95.1000 24.4000 95.4000 24.9000 ;
	    RECT 95.1000 24.0000 95.8000 24.4000 ;
	    RECT 91.9000 23.7000 92.3000 23.8000 ;
	    RECT 93.3000 23.7000 93.7000 23.8000 ;
	    RECT 90.2000 23.1000 90.6000 23.5000 ;
	    RECT 91.9000 23.4000 93.7000 23.7000 ;
	    RECT 93.0000 23.1000 93.3000 23.4000 ;
	    RECT 95.0000 23.1000 95.4000 23.5000 ;
	    RECT 90.2000 22.8000 91.2000 23.1000 ;
	    RECT 90.8000 21.1000 91.2000 22.8000 ;
	    RECT 93.0000 21.1000 93.4000 23.1000 ;
	    RECT 95.1000 21.1000 95.7000 23.1000 ;
	    RECT 97.4000 21.1000 97.8000 25.4000 ;
	    RECT 100.6000 25.4000 101.2000 25.8000 ;
	    RECT 103.0000 25.4000 103.6000 25.8000 ;
	    RECT 104.6000 25.7000 105.0000 27.4000 ;
	    RECT 108.1000 27.1000 108.5000 27.2000 ;
	    RECT 111.0000 27.1000 111.3000 28.2000 ;
	    RECT 113.4000 27.5000 113.8000 29.9000 ;
	    RECT 114.2000 27.8000 114.6000 28.6000 ;
	    RECT 115.0000 28.1000 115.4000 29.9000 ;
	    RECT 116.6000 28.9000 117.0000 29.9000 ;
	    RECT 115.8000 28.1000 116.2000 28.6000 ;
	    RECT 115.0000 27.8000 116.2000 28.1000 ;
	    RECT 112.6000 27.1000 113.4000 27.2000 ;
	    RECT 107.9000 26.8000 113.4000 27.1000 ;
	    RECT 107.0000 26.4000 107.4000 26.5000 ;
	    RECT 105.5000 26.1000 107.4000 26.4000 ;
	    RECT 107.9000 26.2000 108.2000 26.8000 ;
	    RECT 111.5000 26.7000 111.9000 26.8000 ;
	    RECT 111.0000 26.2000 111.4000 26.3000 ;
	    RECT 112.3000 26.2000 112.7000 26.3000 ;
	    RECT 105.5000 26.0000 105.9000 26.1000 ;
	    RECT 107.8000 25.8000 108.2000 26.2000 ;
	    RECT 110.2000 25.9000 112.7000 26.2000 ;
	    RECT 110.2000 25.8000 110.6000 25.9000 ;
	    RECT 106.3000 25.7000 106.7000 25.8000 ;
	    RECT 104.6000 25.4000 106.7000 25.7000 ;
	    RECT 100.6000 25.1000 100.9000 25.4000 ;
	    RECT 103.0000 25.1000 103.3000 25.4000 ;
	    RECT 99.8000 24.8000 100.9000 25.1000 ;
	    RECT 102.2000 24.8000 103.3000 25.1000 ;
	    RECT 99.8000 21.1000 100.2000 24.8000 ;
	    RECT 102.2000 21.1000 102.6000 24.8000 ;
	    RECT 104.6000 21.1000 105.0000 25.4000 ;
	    RECT 107.9000 25.2000 108.2000 25.8000 ;
	    RECT 111.0000 25.5000 113.8000 25.6000 ;
	    RECT 110.9000 25.4000 113.8000 25.5000 ;
	    RECT 107.0000 24.9000 108.2000 25.2000 ;
	    RECT 108.9000 25.3000 113.8000 25.4000 ;
	    RECT 108.9000 25.1000 111.3000 25.3000 ;
	    RECT 107.0000 24.4000 107.3000 24.9000 ;
	    RECT 106.6000 24.0000 107.3000 24.4000 ;
	    RECT 108.1000 24.5000 108.5000 24.6000 ;
	    RECT 108.9000 24.5000 109.2000 25.1000 ;
	    RECT 108.1000 24.2000 109.2000 24.5000 ;
	    RECT 109.5000 24.5000 112.2000 24.8000 ;
	    RECT 109.5000 24.4000 109.9000 24.5000 ;
	    RECT 111.8000 24.4000 112.2000 24.5000 ;
	    RECT 108.7000 23.7000 109.1000 23.8000 ;
	    RECT 110.1000 23.7000 110.5000 23.8000 ;
	    RECT 107.0000 23.1000 107.4000 23.5000 ;
	    RECT 108.7000 23.4000 110.5000 23.7000 ;
	    RECT 109.1000 23.1000 109.4000 23.4000 ;
	    RECT 111.8000 23.1000 112.2000 23.5000 ;
	    RECT 106.7000 21.1000 107.3000 23.1000 ;
	    RECT 109.0000 21.1000 109.4000 23.1000 ;
	    RECT 111.2000 22.8000 112.2000 23.1000 ;
	    RECT 111.2000 21.1000 111.6000 22.8000 ;
	    RECT 113.4000 21.1000 113.8000 25.3000 ;
	    RECT 115.0000 21.1000 115.4000 27.8000 ;
	    RECT 116.7000 27.2000 117.0000 28.9000 ;
	    RECT 118.2000 27.5000 118.6000 29.9000 ;
	    RECT 120.4000 29.2000 120.8000 29.9000 ;
	    RECT 119.8000 28.9000 120.8000 29.2000 ;
	    RECT 122.6000 28.9000 123.0000 29.9000 ;
	    RECT 124.7000 29.2000 125.3000 29.9000 ;
	    RECT 124.6000 28.9000 125.3000 29.2000 ;
	    RECT 119.8000 28.5000 120.2000 28.9000 ;
	    RECT 122.6000 28.6000 122.9000 28.9000 ;
	    RECT 120.6000 28.2000 121.0000 28.6000 ;
	    RECT 121.5000 28.3000 122.9000 28.6000 ;
	    RECT 124.6000 28.5000 125.0000 28.9000 ;
	    RECT 121.5000 28.2000 121.9000 28.3000 ;
	    RECT 115.8000 26.8000 116.2000 27.2000 ;
	    RECT 116.6000 26.8000 117.0000 27.2000 ;
	    RECT 118.6000 27.1000 119.4000 27.2000 ;
	    RECT 120.7000 27.1000 121.0000 28.2000 ;
	    RECT 125.5000 27.7000 125.9000 27.8000 ;
	    RECT 127.0000 27.7000 127.4000 29.9000 ;
	    RECT 125.5000 27.4000 127.4000 27.7000 ;
	    RECT 123.5000 27.1000 123.9000 27.2000 ;
	    RECT 118.6000 26.8000 124.1000 27.1000 ;
	    RECT 115.8000 26.1000 116.1000 26.8000 ;
	    RECT 116.7000 26.1000 117.0000 26.8000 ;
	    RECT 120.1000 26.7000 120.5000 26.8000 ;
	    RECT 119.3000 26.2000 119.7000 26.3000 ;
	    RECT 115.8000 25.8000 117.0000 26.1000 ;
	    RECT 116.7000 25.1000 117.0000 25.8000 ;
	    RECT 117.4000 25.4000 117.8000 26.2000 ;
	    RECT 119.3000 26.1000 121.8000 26.2000 ;
	    RECT 123.0000 26.1000 123.4000 26.2000 ;
	    RECT 119.3000 25.9000 123.4000 26.1000 ;
	    RECT 121.4000 25.8000 123.4000 25.9000 ;
	    RECT 118.2000 25.5000 121.0000 25.6000 ;
	    RECT 118.2000 25.4000 121.1000 25.5000 ;
	    RECT 118.2000 25.3000 123.1000 25.4000 ;
	    RECT 116.6000 24.7000 117.5000 25.1000 ;
	    RECT 117.1000 21.1000 117.5000 24.7000 ;
	    RECT 118.2000 21.1000 118.6000 25.3000 ;
	    RECT 120.7000 25.1000 123.1000 25.3000 ;
	    RECT 119.8000 24.5000 122.5000 24.8000 ;
	    RECT 119.8000 24.4000 120.2000 24.5000 ;
	    RECT 122.1000 24.4000 122.5000 24.5000 ;
	    RECT 122.8000 24.5000 123.1000 25.1000 ;
	    RECT 123.8000 25.2000 124.1000 26.8000 ;
	    RECT 124.6000 26.4000 125.0000 26.5000 ;
	    RECT 124.6000 26.1000 126.5000 26.4000 ;
	    RECT 126.1000 26.0000 126.5000 26.1000 ;
	    RECT 125.3000 25.7000 125.7000 25.8000 ;
	    RECT 127.0000 25.7000 127.4000 27.4000 ;
	    RECT 128.6000 28.8000 129.0000 29.9000 ;
	    RECT 128.6000 27.2000 128.9000 28.8000 ;
	    RECT 129.4000 27.8000 129.8000 28.6000 ;
	    RECT 131.8000 27.9000 132.2000 29.9000 ;
	    RECT 134.2000 28.9000 134.6000 29.9000 ;
	    RECT 132.5000 28.2000 132.9000 28.6000 ;
	    RECT 132.6000 28.1000 133.0000 28.2000 ;
	    RECT 134.2000 28.1000 134.5000 28.9000 ;
	    RECT 128.6000 26.8000 129.0000 27.2000 ;
	    RECT 125.3000 25.4000 127.4000 25.7000 ;
	    RECT 127.8000 25.4000 128.2000 26.2000 ;
	    RECT 123.8000 24.9000 125.0000 25.2000 ;
	    RECT 123.5000 24.5000 123.9000 24.6000 ;
	    RECT 122.8000 24.2000 123.9000 24.5000 ;
	    RECT 124.7000 24.4000 125.0000 24.9000 ;
	    RECT 124.7000 24.0000 125.4000 24.4000 ;
	    RECT 121.5000 23.7000 121.9000 23.8000 ;
	    RECT 122.9000 23.7000 123.3000 23.8000 ;
	    RECT 119.8000 23.1000 120.2000 23.5000 ;
	    RECT 121.5000 23.4000 123.3000 23.7000 ;
	    RECT 122.6000 23.1000 122.9000 23.4000 ;
	    RECT 124.6000 23.1000 125.0000 23.5000 ;
	    RECT 119.8000 22.8000 120.8000 23.1000 ;
	    RECT 120.4000 21.1000 120.8000 22.8000 ;
	    RECT 122.6000 21.1000 123.0000 23.1000 ;
	    RECT 124.7000 21.1000 125.3000 23.1000 ;
	    RECT 127.0000 21.1000 127.4000 25.4000 ;
	    RECT 128.6000 25.1000 128.9000 26.8000 ;
	    RECT 131.0000 26.4000 131.4000 27.2000 ;
	    RECT 130.2000 26.1000 130.6000 26.2000 ;
	    RECT 131.8000 26.1000 132.1000 27.9000 ;
	    RECT 132.6000 27.8000 134.5000 28.1000 ;
	    RECT 135.0000 27.8000 135.4000 28.6000 ;
	    RECT 134.2000 27.2000 134.5000 27.8000 ;
	    RECT 135.8000 27.5000 136.2000 29.9000 ;
	    RECT 138.0000 29.2000 138.4000 29.9000 ;
	    RECT 137.4000 28.9000 138.4000 29.2000 ;
	    RECT 140.2000 28.9000 140.6000 29.9000 ;
	    RECT 142.3000 29.2000 142.9000 29.9000 ;
	    RECT 142.2000 28.9000 142.9000 29.2000 ;
	    RECT 137.4000 28.5000 137.8000 28.9000 ;
	    RECT 140.2000 28.6000 140.5000 28.9000 ;
	    RECT 138.2000 28.2000 138.6000 28.6000 ;
	    RECT 139.1000 28.3000 140.5000 28.6000 ;
	    RECT 142.2000 28.5000 142.6000 28.9000 ;
	    RECT 139.1000 28.2000 139.5000 28.3000 ;
	    RECT 138.3000 27.2000 138.6000 28.2000 ;
	    RECT 143.1000 27.7000 143.5000 27.8000 ;
	    RECT 144.6000 27.7000 145.0000 29.9000 ;
	    RECT 143.1000 27.4000 145.0000 27.7000 ;
	    RECT 134.2000 26.8000 134.6000 27.2000 ;
	    RECT 136.2000 27.1000 137.0000 27.2000 ;
	    RECT 138.2000 27.1000 138.6000 27.2000 ;
	    RECT 141.1000 27.1000 141.5000 27.2000 ;
	    RECT 136.2000 26.8000 141.7000 27.1000 ;
	    RECT 132.6000 26.1000 133.0000 26.2000 ;
	    RECT 130.2000 25.8000 131.0000 26.1000 ;
	    RECT 131.8000 25.8000 133.0000 26.1000 ;
	    RECT 130.6000 25.6000 131.0000 25.8000 ;
	    RECT 132.6000 25.1000 132.9000 25.8000 ;
	    RECT 133.4000 25.4000 133.8000 26.2000 ;
	    RECT 134.2000 25.1000 134.5000 26.8000 ;
	    RECT 137.7000 26.7000 138.1000 26.8000 ;
	    RECT 136.9000 26.2000 137.3000 26.3000 ;
	    RECT 136.9000 25.9000 139.4000 26.2000 ;
	    RECT 139.0000 25.8000 139.4000 25.9000 ;
	    RECT 135.8000 25.5000 138.6000 25.6000 ;
	    RECT 135.8000 25.4000 138.7000 25.5000 ;
	    RECT 135.8000 25.3000 140.7000 25.4000 ;
	    RECT 128.1000 24.7000 129.0000 25.1000 ;
	    RECT 130.2000 24.8000 132.2000 25.1000 ;
	    RECT 128.1000 21.1000 128.5000 24.7000 ;
	    RECT 130.2000 21.1000 130.6000 24.8000 ;
	    RECT 131.8000 21.1000 132.2000 24.8000 ;
	    RECT 132.6000 21.1000 133.0000 25.1000 ;
	    RECT 133.7000 24.7000 134.6000 25.1000 ;
	    RECT 133.7000 21.1000 134.1000 24.7000 ;
	    RECT 135.8000 21.1000 136.2000 25.3000 ;
	    RECT 138.3000 25.1000 140.7000 25.3000 ;
	    RECT 137.4000 24.5000 140.1000 24.8000 ;
	    RECT 137.4000 24.4000 137.8000 24.5000 ;
	    RECT 139.7000 24.4000 140.1000 24.5000 ;
	    RECT 140.4000 24.5000 140.7000 25.1000 ;
	    RECT 141.4000 25.2000 141.7000 26.8000 ;
	    RECT 142.2000 26.4000 142.6000 26.5000 ;
	    RECT 142.2000 26.1000 144.1000 26.4000 ;
	    RECT 143.7000 26.0000 144.1000 26.1000 ;
	    RECT 142.9000 25.7000 143.3000 25.8000 ;
	    RECT 144.6000 25.7000 145.0000 27.4000 ;
	    RECT 145.4000 27.6000 145.8000 29.9000 ;
	    RECT 145.4000 27.3000 146.5000 27.6000 ;
	    RECT 145.4000 25.8000 145.8000 26.6000 ;
	    RECT 146.2000 25.8000 146.5000 27.3000 ;
	    RECT 142.9000 25.4000 145.0000 25.7000 ;
	    RECT 141.4000 24.9000 142.6000 25.2000 ;
	    RECT 141.1000 24.5000 141.5000 24.6000 ;
	    RECT 140.4000 24.2000 141.5000 24.5000 ;
	    RECT 142.3000 24.4000 142.6000 24.9000 ;
	    RECT 142.3000 24.0000 143.0000 24.4000 ;
	    RECT 139.1000 23.7000 139.5000 23.8000 ;
	    RECT 140.5000 23.7000 140.9000 23.8000 ;
	    RECT 137.4000 23.1000 137.8000 23.5000 ;
	    RECT 139.1000 23.4000 140.9000 23.7000 ;
	    RECT 140.2000 23.1000 140.5000 23.4000 ;
	    RECT 142.2000 23.1000 142.6000 23.5000 ;
	    RECT 137.4000 22.8000 138.4000 23.1000 ;
	    RECT 138.0000 21.1000 138.4000 22.8000 ;
	    RECT 140.2000 21.1000 140.6000 23.1000 ;
	    RECT 142.3000 21.1000 142.9000 23.1000 ;
	    RECT 144.6000 21.1000 145.0000 25.4000 ;
	    RECT 146.2000 25.4000 146.8000 25.8000 ;
	    RECT 146.2000 25.1000 146.5000 25.4000 ;
	    RECT 145.4000 24.8000 146.5000 25.1000 ;
	    RECT 145.4000 21.1000 145.8000 24.8000 ;
	    RECT 0.6000 15.6000 1.0000 19.9000 ;
	    RECT 2.7000 17.9000 3.3000 19.9000 ;
	    RECT 5.0000 17.9000 5.4000 19.9000 ;
	    RECT 7.2000 18.2000 7.6000 19.9000 ;
	    RECT 7.2000 17.9000 8.2000 18.2000 ;
	    RECT 3.0000 17.5000 3.4000 17.9000 ;
	    RECT 5.1000 17.6000 5.4000 17.9000 ;
	    RECT 4.7000 17.3000 6.5000 17.6000 ;
	    RECT 7.8000 17.5000 8.2000 17.9000 ;
	    RECT 4.7000 17.2000 5.1000 17.3000 ;
	    RECT 6.1000 17.2000 6.5000 17.3000 ;
	    RECT 2.6000 16.6000 3.3000 17.0000 ;
	    RECT 3.0000 16.1000 3.3000 16.6000 ;
	    RECT 4.1000 16.5000 5.2000 16.8000 ;
	    RECT 4.1000 16.4000 4.5000 16.5000 ;
	    RECT 3.0000 15.8000 4.2000 16.1000 ;
	    RECT 0.6000 15.3000 2.7000 15.6000 ;
	    RECT 0.6000 13.6000 1.0000 15.3000 ;
	    RECT 2.3000 15.2000 2.7000 15.3000 ;
	    RECT 1.5000 14.9000 1.9000 15.0000 ;
	    RECT 1.5000 14.6000 3.4000 14.9000 ;
	    RECT 3.0000 14.5000 3.4000 14.6000 ;
	    RECT 3.9000 14.2000 4.2000 15.8000 ;
	    RECT 4.9000 15.9000 5.2000 16.5000 ;
	    RECT 5.5000 16.5000 5.9000 16.6000 ;
	    RECT 7.8000 16.5000 8.2000 16.6000 ;
	    RECT 5.5000 16.2000 8.2000 16.5000 ;
	    RECT 4.9000 15.7000 7.3000 15.9000 ;
	    RECT 9.4000 15.7000 9.8000 19.9000 ;
	    RECT 4.9000 15.6000 9.8000 15.7000 ;
	    RECT 6.9000 15.5000 9.8000 15.6000 ;
	    RECT 7.0000 15.4000 9.8000 15.5000 ;
	    RECT 10.2000 15.6000 10.6000 19.9000 ;
	    RECT 12.3000 17.9000 12.9000 19.9000 ;
	    RECT 14.6000 17.9000 15.0000 19.9000 ;
	    RECT 16.8000 18.2000 17.2000 19.9000 ;
	    RECT 16.8000 17.9000 17.8000 18.2000 ;
	    RECT 12.6000 17.5000 13.0000 17.9000 ;
	    RECT 14.7000 17.6000 15.0000 17.9000 ;
	    RECT 14.3000 17.3000 16.1000 17.6000 ;
	    RECT 17.4000 17.5000 17.8000 17.9000 ;
	    RECT 14.3000 17.2000 14.7000 17.3000 ;
	    RECT 15.7000 17.2000 16.1000 17.3000 ;
	    RECT 12.2000 16.6000 12.9000 17.0000 ;
	    RECT 12.6000 16.1000 12.9000 16.6000 ;
	    RECT 13.7000 16.5000 14.8000 16.8000 ;
	    RECT 13.7000 16.4000 14.1000 16.5000 ;
	    RECT 12.6000 15.8000 13.8000 16.1000 ;
	    RECT 10.2000 15.3000 12.3000 15.6000 ;
	    RECT 7.5000 14.2000 7.9000 14.3000 ;
	    RECT 3.9000 13.9000 9.4000 14.2000 ;
	    RECT 4.1000 13.8000 4.5000 13.9000 ;
	    RECT 0.6000 13.3000 2.5000 13.6000 ;
	    RECT 0.6000 11.1000 1.0000 13.3000 ;
	    RECT 2.1000 13.2000 2.5000 13.3000 ;
	    RECT 7.0000 12.8000 7.3000 13.9000 ;
	    RECT 8.6000 13.8000 9.4000 13.9000 ;
	    RECT 10.2000 13.6000 10.6000 15.3000 ;
	    RECT 11.9000 15.2000 12.3000 15.3000 ;
	    RECT 13.5000 15.2000 13.8000 15.8000 ;
	    RECT 14.5000 15.9000 14.8000 16.5000 ;
	    RECT 15.1000 16.5000 15.5000 16.6000 ;
	    RECT 17.4000 16.5000 17.8000 16.6000 ;
	    RECT 15.1000 16.2000 17.8000 16.5000 ;
	    RECT 14.5000 15.7000 16.9000 15.9000 ;
	    RECT 19.0000 15.7000 19.4000 19.9000 ;
	    RECT 19.8000 17.9000 20.2000 19.9000 ;
	    RECT 19.9000 17.8000 20.2000 17.9000 ;
	    RECT 21.4000 17.9000 21.8000 19.9000 ;
	    RECT 21.4000 17.8000 21.7000 17.9000 ;
	    RECT 19.9000 17.5000 21.7000 17.8000 ;
	    RECT 19.9000 16.2000 20.2000 17.5000 ;
	    RECT 20.6000 16.4000 21.0000 17.2000 ;
	    RECT 19.8000 15.8000 20.2000 16.2000 ;
	    RECT 14.5000 15.6000 19.4000 15.7000 ;
	    RECT 16.5000 15.5000 19.4000 15.6000 ;
	    RECT 16.6000 15.4000 19.4000 15.5000 ;
	    RECT 19.9000 15.2000 20.2000 15.8000 ;
	    RECT 22.2000 15.4000 22.6000 16.2000 ;
	    RECT 11.1000 14.9000 11.5000 15.0000 ;
	    RECT 11.1000 14.6000 13.0000 14.9000 ;
	    RECT 13.4000 14.8000 13.8000 15.2000 ;
	    RECT 15.8000 15.1000 16.2000 15.2000 ;
	    RECT 15.8000 14.8000 18.3000 15.1000 ;
	    RECT 19.8000 14.8000 20.2000 15.2000 ;
	    RECT 21.0000 14.8000 21.8000 15.2000 ;
	    RECT 12.6000 14.5000 13.0000 14.6000 ;
	    RECT 13.5000 14.2000 13.8000 14.8000 ;
	    RECT 16.6000 14.7000 17.0000 14.8000 ;
	    RECT 17.9000 14.7000 18.3000 14.8000 ;
	    RECT 17.1000 14.2000 17.5000 14.3000 ;
	    RECT 19.9000 14.2000 20.2000 14.8000 ;
	    RECT 13.5000 13.9000 19.0000 14.2000 ;
	    RECT 19.9000 14.1000 20.7000 14.2000 ;
	    RECT 19.9000 13.9000 20.8000 14.1000 ;
	    RECT 13.7000 13.8000 14.1000 13.9000 ;
	    RECT 6.1000 12.7000 6.5000 12.8000 ;
	    RECT 3.0000 12.1000 3.4000 12.5000 ;
	    RECT 5.1000 12.4000 6.5000 12.7000 ;
	    RECT 7.0000 12.4000 7.4000 12.8000 ;
	    RECT 5.1000 12.1000 5.4000 12.4000 ;
	    RECT 7.8000 12.1000 8.2000 12.5000 ;
	    RECT 2.7000 11.8000 3.4000 12.1000 ;
	    RECT 2.7000 11.1000 3.3000 11.8000 ;
	    RECT 5.0000 11.1000 5.4000 12.1000 ;
	    RECT 7.2000 11.8000 8.2000 12.1000 ;
	    RECT 7.2000 11.1000 7.6000 11.8000 ;
	    RECT 9.4000 11.1000 9.8000 13.5000 ;
	    RECT 10.2000 13.3000 12.1000 13.6000 ;
	    RECT 10.2000 11.1000 10.6000 13.3000 ;
	    RECT 11.7000 13.2000 12.1000 13.3000 ;
	    RECT 16.6000 12.8000 16.9000 13.9000 ;
	    RECT 18.2000 13.8000 19.0000 13.9000 ;
	    RECT 15.7000 12.7000 16.1000 12.8000 ;
	    RECT 12.6000 12.1000 13.0000 12.5000 ;
	    RECT 14.7000 12.4000 16.1000 12.7000 ;
	    RECT 16.6000 12.4000 17.0000 12.8000 ;
	    RECT 14.7000 12.1000 15.0000 12.4000 ;
	    RECT 17.4000 12.1000 17.8000 12.5000 ;
	    RECT 12.3000 11.8000 13.0000 12.1000 ;
	    RECT 12.3000 11.1000 12.9000 11.8000 ;
	    RECT 14.6000 11.1000 15.0000 12.1000 ;
	    RECT 16.8000 11.8000 17.8000 12.1000 ;
	    RECT 16.8000 11.1000 17.2000 11.8000 ;
	    RECT 19.0000 11.1000 19.4000 13.5000 ;
	    RECT 20.4000 11.1000 20.8000 13.9000 ;
	    RECT 23.0000 11.1000 23.4000 19.9000 ;
	    RECT 25.4000 17.9000 25.8000 19.9000 ;
	    RECT 25.5000 17.8000 25.8000 17.9000 ;
	    RECT 27.0000 17.9000 27.4000 19.9000 ;
	    RECT 27.0000 17.8000 27.3000 17.9000 ;
	    RECT 25.5000 17.5000 27.3000 17.8000 ;
	    RECT 26.2000 16.4000 26.6000 17.2000 ;
	    RECT 27.0000 16.2000 27.3000 17.5000 ;
	    RECT 29.1000 16.3000 29.5000 19.9000 ;
	    RECT 27.0000 15.8000 27.4000 16.2000 ;
	    RECT 28.6000 15.9000 29.5000 16.3000 ;
	    RECT 28.6000 15.8000 29.0000 15.9000 ;
	    RECT 25.4000 14.8000 26.2000 15.2000 ;
	    RECT 27.0000 14.2000 27.3000 15.8000 ;
	    RECT 28.7000 14.2000 29.0000 15.8000 ;
	    RECT 29.4000 14.8000 29.8000 15.6000 ;
	    RECT 26.5000 14.1000 27.3000 14.2000 ;
	    RECT 26.4000 13.9000 27.3000 14.1000 ;
	    RECT 23.8000 12.4000 24.2000 13.2000 ;
	    RECT 26.4000 11.1000 26.8000 13.9000 ;
	    RECT 28.6000 13.8000 29.0000 14.2000 ;
	    RECT 27.8000 12.4000 28.2000 13.2000 ;
	    RECT 28.7000 12.1000 29.0000 13.8000 ;
	    RECT 30.2000 13.4000 30.6000 14.2000 ;
	    RECT 31.0000 13.1000 31.4000 19.9000 ;
	    RECT 33.0000 16.8000 33.4000 17.2000 ;
	    RECT 31.8000 15.8000 32.2000 16.6000 ;
	    RECT 33.0000 16.2000 33.3000 16.8000 ;
	    RECT 33.7000 16.2000 34.1000 19.9000 ;
	    RECT 37.1000 16.3000 37.5000 19.9000 ;
	    RECT 32.6000 15.9000 33.3000 16.2000 ;
	    RECT 33.6000 15.9000 34.1000 16.2000 ;
	    RECT 36.6000 15.9000 37.5000 16.3000 ;
	    RECT 32.6000 15.8000 33.0000 15.9000 ;
	    RECT 31.8000 14.8000 32.2000 15.2000 ;
	    RECT 31.8000 14.1000 32.1000 14.8000 ;
	    RECT 33.6000 14.2000 33.9000 15.9000 ;
	    RECT 34.2000 15.1000 34.6000 15.2000 ;
	    RECT 35.8000 15.1000 36.2000 15.2000 ;
	    RECT 34.2000 14.8000 36.2000 15.1000 ;
	    RECT 34.2000 14.4000 34.6000 14.8000 ;
	    RECT 36.7000 14.2000 37.0000 15.9000 ;
	    RECT 32.6000 14.1000 33.9000 14.2000 ;
	    RECT 35.0000 14.1000 35.4000 14.2000 ;
	    RECT 31.8000 13.8000 33.9000 14.1000 ;
	    RECT 34.6000 13.8000 35.4000 14.1000 ;
	    RECT 36.6000 13.8000 37.0000 14.2000 ;
	    RECT 37.4000 15.1000 37.8000 15.6000 ;
	    RECT 38.2000 15.1000 38.6000 19.9000 ;
	    RECT 37.4000 14.8000 38.6000 15.1000 ;
	    RECT 37.4000 14.2000 37.7000 14.8000 ;
	    RECT 37.4000 13.8000 37.8000 14.2000 ;
	    RECT 32.7000 13.1000 33.0000 13.8000 ;
	    RECT 34.6000 13.6000 35.0000 13.8000 ;
	    RECT 33.5000 13.1000 35.3000 13.3000 ;
	    RECT 31.0000 12.8000 31.9000 13.1000 ;
	    RECT 28.6000 11.1000 29.0000 12.1000 ;
	    RECT 31.5000 11.1000 31.9000 12.8000 ;
	    RECT 32.6000 11.1000 33.0000 13.1000 ;
	    RECT 33.4000 13.0000 35.4000 13.1000 ;
	    RECT 33.4000 11.1000 33.8000 13.0000 ;
	    RECT 35.0000 11.1000 35.4000 13.0000 ;
	    RECT 35.8000 12.4000 36.2000 13.2000 ;
	    RECT 36.7000 12.2000 37.0000 13.8000 ;
	    RECT 36.6000 11.1000 37.0000 12.2000 ;
	    RECT 38.2000 11.1000 38.6000 14.8000 ;
	    RECT 39.0000 13.1000 39.4000 13.2000 ;
	    RECT 40.6000 13.1000 41.0000 19.9000 ;
	    RECT 43.0000 17.9000 43.4000 19.9000 ;
	    RECT 43.1000 17.8000 43.4000 17.9000 ;
	    RECT 44.6000 17.9000 45.0000 19.9000 ;
	    RECT 44.6000 17.8000 44.9000 17.9000 ;
	    RECT 43.1000 17.5000 44.9000 17.8000 ;
	    RECT 44.6000 16.2000 44.9000 17.5000 ;
	    RECT 45.7000 16.3000 46.1000 19.9000 ;
	    RECT 44.6000 15.8000 45.0000 16.2000 ;
	    RECT 45.7000 15.9000 46.6000 16.3000 ;
	    RECT 50.7000 15.9000 51.7000 19.9000 ;
	    RECT 54.5000 19.2000 54.9000 19.9000 ;
	    RECT 54.5000 18.8000 55.4000 19.2000 ;
	    RECT 53.8000 16.8000 54.2000 17.2000 ;
	    RECT 53.8000 16.2000 54.1000 16.8000 ;
	    RECT 54.5000 16.2000 54.9000 18.8000 ;
	    RECT 53.4000 15.9000 54.1000 16.2000 ;
	    RECT 54.4000 15.9000 54.9000 16.2000 ;
	    RECT 44.6000 14.2000 44.9000 15.8000 ;
	    RECT 46.2000 15.1000 46.5000 15.9000 ;
	    RECT 50.2000 15.1000 50.6000 15.2000 ;
	    RECT 46.2000 14.8000 50.6000 15.1000 ;
	    RECT 46.2000 14.2000 46.5000 14.8000 ;
	    RECT 50.2000 14.4000 50.6000 14.8000 ;
	    RECT 51.0000 14.2000 51.3000 15.9000 ;
	    RECT 53.4000 15.8000 53.8000 15.9000 ;
	    RECT 51.8000 14.4000 52.2000 15.2000 ;
	    RECT 44.1000 14.1000 44.9000 14.2000 ;
	    RECT 39.0000 12.8000 41.0000 13.1000 ;
	    RECT 44.0000 13.9000 44.9000 14.1000 ;
	    RECT 39.0000 12.4000 39.4000 12.8000 ;
	    RECT 40.1000 11.1000 40.5000 12.8000 ;
	    RECT 44.0000 12.2000 44.4000 13.9000 ;
	    RECT 45.4000 13.8000 45.8000 14.2000 ;
	    RECT 46.2000 13.8000 46.6000 14.2000 ;
	    RECT 49.4000 14.1000 49.8000 14.2000 ;
	    RECT 51.0000 14.1000 51.4000 14.2000 ;
	    RECT 49.4000 13.8000 50.2000 14.1000 ;
	    RECT 51.0000 13.8000 52.2000 14.1000 ;
	    RECT 52.6000 13.8000 53.0000 14.6000 ;
	    RECT 54.4000 14.2000 54.7000 15.9000 ;
	    RECT 57.4000 15.1000 57.8000 19.9000 ;
	    RECT 58.2000 16.2000 58.6000 19.9000 ;
	    RECT 59.8000 16.2000 60.2000 19.9000 ;
	    RECT 58.2000 15.9000 60.2000 16.2000 ;
	    RECT 60.6000 15.9000 61.0000 19.9000 ;
	    RECT 61.7000 19.2000 62.1000 19.9000 ;
	    RECT 61.4000 18.8000 62.1000 19.2000 ;
	    RECT 61.7000 16.3000 62.1000 18.8000 ;
	    RECT 61.7000 15.9000 62.6000 16.3000 ;
	    RECT 58.6000 15.2000 59.0000 15.4000 ;
	    RECT 60.6000 15.2000 60.9000 15.9000 ;
	    RECT 58.2000 15.1000 59.0000 15.2000 ;
	    RECT 57.4000 14.9000 59.0000 15.1000 ;
	    RECT 59.8000 15.1000 61.0000 15.2000 ;
	    RECT 61.4000 15.1000 61.8000 15.6000 ;
	    RECT 59.8000 14.9000 61.8000 15.1000 ;
	    RECT 57.4000 14.8000 58.6000 14.9000 ;
	    RECT 53.4000 13.8000 54.7000 14.2000 ;
	    RECT 55.8000 14.1000 56.2000 14.2000 ;
	    RECT 55.4000 13.8000 56.2000 14.1000 ;
	    RECT 45.4000 13.1000 45.7000 13.8000 ;
	    RECT 46.2000 13.1000 46.5000 13.8000 ;
	    RECT 49.8000 13.6000 50.2000 13.8000 ;
	    RECT 49.5000 13.1000 51.3000 13.3000 ;
	    RECT 51.9000 13.2000 52.2000 13.8000 ;
	    RECT 45.4000 12.8000 46.5000 13.1000 ;
	    RECT 43.8000 11.8000 44.4000 12.2000 ;
	    RECT 44.0000 11.1000 44.4000 11.8000 ;
	    RECT 46.2000 12.1000 46.5000 12.8000 ;
	    RECT 49.4000 13.0000 51.4000 13.1000 ;
	    RECT 46.2000 11.1000 46.6000 12.1000 ;
	    RECT 49.4000 11.1000 49.8000 13.0000 ;
	    RECT 51.0000 11.4000 51.4000 13.0000 ;
	    RECT 51.8000 11.7000 52.2000 13.2000 ;
	    RECT 53.5000 13.1000 53.8000 13.8000 ;
	    RECT 55.4000 13.6000 55.8000 13.8000 ;
	    RECT 54.3000 13.1000 56.1000 13.3000 ;
	    RECT 52.6000 11.4000 53.0000 13.1000 ;
	    RECT 51.0000 11.1000 53.0000 11.4000 ;
	    RECT 53.4000 11.1000 53.8000 13.1000 ;
	    RECT 54.2000 13.0000 56.2000 13.1000 ;
	    RECT 54.2000 11.1000 54.6000 13.0000 ;
	    RECT 55.8000 11.1000 56.2000 13.0000 ;
	    RECT 57.4000 11.1000 57.8000 14.8000 ;
	    RECT 59.0000 13.8000 59.4000 14.6000 ;
	    RECT 59.8000 13.1000 60.1000 14.9000 ;
	    RECT 60.6000 14.8000 61.8000 14.9000 ;
	    RECT 62.2000 14.2000 62.5000 15.9000 ;
	    RECT 62.2000 13.8000 62.6000 14.2000 ;
	    RECT 59.8000 11.1000 60.2000 13.1000 ;
	    RECT 60.6000 12.8000 61.0000 13.2000 ;
	    RECT 60.5000 12.4000 60.9000 12.8000 ;
	    RECT 62.2000 12.1000 62.5000 13.8000 ;
	    RECT 63.8000 13.4000 64.2000 14.2000 ;
	    RECT 63.0000 12.4000 63.4000 13.2000 ;
	    RECT 64.6000 13.1000 65.0000 19.9000 ;
	    RECT 65.4000 15.8000 65.8000 16.6000 ;
	    RECT 66.5000 16.3000 66.9000 19.9000 ;
	    RECT 66.5000 15.9000 67.4000 16.3000 ;
	    RECT 69.4000 16.1000 69.8000 19.9000 ;
	    RECT 70.2000 16.1000 70.6000 16.6000 ;
	    RECT 66.2000 14.8000 66.6000 15.6000 ;
	    RECT 67.0000 14.2000 67.3000 15.9000 ;
	    RECT 69.4000 15.8000 70.6000 16.1000 ;
	    RECT 68.6000 14.8000 69.0000 15.2000 ;
	    RECT 67.0000 14.1000 67.4000 14.2000 ;
	    RECT 68.6000 14.1000 68.9000 14.8000 ;
	    RECT 67.0000 13.8000 68.9000 14.1000 ;
	    RECT 64.6000 12.8000 65.5000 13.1000 ;
	    RECT 62.2000 11.1000 62.6000 12.1000 ;
	    RECT 65.1000 11.1000 65.5000 12.8000 ;
	    RECT 67.0000 12.1000 67.3000 13.8000 ;
	    RECT 67.0000 11.1000 67.4000 12.1000 ;
	    RECT 69.4000 11.1000 69.8000 15.8000 ;
	    RECT 71.0000 13.1000 71.4000 19.9000 ;
	    RECT 72.6000 16.9000 73.0000 19.9000 ;
	    RECT 72.7000 16.6000 73.0000 16.9000 ;
	    RECT 74.2000 19.6000 76.2000 19.9000 ;
	    RECT 74.2000 16.9000 74.6000 19.6000 ;
	    RECT 75.0000 16.9000 75.4000 19.3000 ;
	    RECT 75.8000 17.0000 76.2000 19.6000 ;
	    RECT 76.7000 19.6000 78.5000 19.9000 ;
	    RECT 76.7000 19.5000 77.0000 19.6000 ;
	    RECT 74.2000 16.6000 74.5000 16.9000 ;
	    RECT 72.7000 16.3000 74.5000 16.6000 ;
	    RECT 75.1000 16.7000 75.4000 16.9000 ;
	    RECT 76.6000 16.7000 77.0000 19.5000 ;
	    RECT 78.2000 19.5000 78.5000 19.6000 ;
	    RECT 75.1000 16.5000 77.0000 16.7000 ;
	    RECT 77.4000 16.5000 77.8000 19.3000 ;
	    RECT 78.2000 16.5000 78.6000 19.5000 ;
	    RECT 79.0000 16.9000 79.4000 19.9000 ;
	    RECT 79.1000 16.6000 79.4000 16.9000 ;
	    RECT 80.6000 19.6000 82.6000 19.9000 ;
	    RECT 80.6000 16.9000 81.0000 19.6000 ;
	    RECT 81.4000 16.9000 81.8000 19.3000 ;
	    RECT 82.2000 17.0000 82.6000 19.6000 ;
	    RECT 83.1000 19.6000 84.9000 19.9000 ;
	    RECT 83.1000 19.5000 83.4000 19.6000 ;
	    RECT 80.6000 16.6000 80.9000 16.9000 ;
	    RECT 75.1000 16.4000 76.9000 16.5000 ;
	    RECT 77.4000 16.2000 77.7000 16.5000 ;
	    RECT 79.1000 16.3000 80.9000 16.6000 ;
	    RECT 81.5000 16.7000 81.8000 16.9000 ;
	    RECT 83.0000 16.7000 83.4000 19.5000 ;
	    RECT 84.6000 19.5000 84.9000 19.6000 ;
	    RECT 81.5000 16.5000 83.4000 16.7000 ;
	    RECT 83.8000 16.5000 84.2000 19.3000 ;
	    RECT 84.6000 16.5000 85.0000 19.5000 ;
	    RECT 85.4000 16.9000 85.8000 19.9000 ;
	    RECT 85.5000 16.6000 85.8000 16.9000 ;
	    RECT 87.0000 19.6000 89.0000 19.9000 ;
	    RECT 87.0000 16.9000 87.4000 19.6000 ;
	    RECT 87.8000 16.9000 88.2000 19.3000 ;
	    RECT 88.6000 17.0000 89.0000 19.6000 ;
	    RECT 89.5000 19.6000 91.3000 19.9000 ;
	    RECT 89.5000 19.5000 89.8000 19.6000 ;
	    RECT 87.0000 16.6000 87.3000 16.9000 ;
	    RECT 81.5000 16.4000 83.3000 16.5000 ;
	    RECT 83.8000 16.2000 84.1000 16.5000 ;
	    RECT 85.5000 16.3000 87.3000 16.6000 ;
	    RECT 87.9000 16.7000 88.2000 16.9000 ;
	    RECT 89.4000 16.7000 89.8000 19.5000 ;
	    RECT 91.0000 19.5000 91.3000 19.6000 ;
	    RECT 87.9000 16.5000 89.8000 16.7000 ;
	    RECT 90.2000 16.5000 90.6000 19.3000 ;
	    RECT 91.0000 16.5000 91.4000 19.5000 ;
	    RECT 87.9000 16.4000 89.7000 16.5000 ;
	    RECT 90.2000 16.2000 90.5000 16.5000 ;
	    RECT 92.1000 16.3000 92.5000 19.9000 ;
	    RECT 94.5000 16.3000 94.9000 19.9000 ;
	    RECT 77.4000 16.1000 77.8000 16.2000 ;
	    RECT 83.8000 16.1000 84.2000 16.2000 ;
	    RECT 90.2000 16.1000 90.6000 16.2000 ;
	    RECT 76.1000 15.8000 77.8000 16.1000 ;
	    RECT 82.5000 15.8000 84.2000 16.1000 ;
	    RECT 88.9000 15.8000 90.6000 16.1000 ;
	    RECT 92.1000 15.9000 93.0000 16.3000 ;
	    RECT 94.5000 15.9000 95.4000 16.3000 ;
	    RECT 72.6000 15.1000 73.0000 15.2000 ;
	    RECT 75.0000 15.1000 75.8000 15.2000 ;
	    RECT 72.6000 14.8000 75.8000 15.1000 ;
	    RECT 74.2000 13.8000 75.0000 14.2000 ;
	    RECT 70.5000 12.8000 71.4000 13.1000 ;
	    RECT 73.4000 13.1000 74.3000 13.2000 ;
	    RECT 75.0000 13.1000 75.4000 13.2000 ;
	    RECT 73.4000 12.8000 75.4000 13.1000 ;
	    RECT 70.5000 11.1000 70.9000 12.8000 ;
	    RECT 76.1000 12.5000 76.4000 15.8000 ;
	    RECT 77.4000 15.1000 77.8000 15.2000 ;
	    RECT 81.4000 15.1000 82.2000 15.2000 ;
	    RECT 77.4000 14.8000 82.2000 15.1000 ;
	    RECT 80.6000 13.8000 81.4000 14.2000 ;
	    RECT 79.0000 13.1000 79.4000 13.2000 ;
	    RECT 79.8000 13.1000 80.7000 13.2000 ;
	    RECT 79.0000 12.8000 80.7000 13.1000 ;
	    RECT 82.5000 12.5000 82.8000 15.8000 ;
	    RECT 87.8000 14.8000 88.6000 15.2000 ;
	    RECT 84.6000 14.1000 85.0000 14.2000 ;
	    RECT 87.0000 14.1000 87.8000 14.2000 ;
	    RECT 84.6000 13.8000 87.8000 14.1000 ;
	    RECT 85.4000 13.1000 85.8000 13.2000 ;
	    RECT 86.2000 13.1000 87.1000 13.2000 ;
	    RECT 85.4000 12.8000 87.1000 13.1000 ;
	    RECT 88.9000 12.5000 89.2000 15.8000 ;
	    RECT 91.0000 15.1000 91.4000 15.2000 ;
	    RECT 91.8000 15.1000 92.2000 15.6000 ;
	    RECT 91.0000 14.8000 92.2000 15.1000 ;
	    RECT 74.4000 12.2000 76.4000 12.5000 ;
	    RECT 80.8000 12.2000 82.8000 12.5000 ;
	    RECT 87.2000 12.2000 89.2000 12.5000 ;
	    RECT 74.2000 11.8000 74.7000 12.2000 ;
	    RECT 75.8000 12.1000 76.4000 12.2000 ;
	    RECT 74.2000 11.1000 74.6000 11.8000 ;
	    RECT 75.8000 11.1000 76.2000 12.1000 ;
	    RECT 80.6000 11.8000 81.1000 12.2000 ;
	    RECT 82.2000 12.1000 82.8000 12.2000 ;
	    RECT 80.6000 11.1000 81.0000 11.8000 ;
	    RECT 82.2000 11.1000 82.6000 12.1000 ;
	    RECT 87.0000 11.8000 87.5000 12.2000 ;
	    RECT 88.6000 12.1000 89.2000 12.2000 ;
	    RECT 92.6000 14.2000 92.9000 15.9000 ;
	    RECT 94.2000 14.8000 94.6000 15.6000 ;
	    RECT 95.0000 14.2000 95.3000 15.9000 ;
	    RECT 96.6000 15.8000 97.0000 16.6000 ;
	    RECT 92.6000 13.8000 93.0000 14.2000 ;
	    RECT 95.0000 13.8000 95.4000 14.2000 ;
	    RECT 95.8000 13.8000 96.2000 14.2000 ;
	    RECT 92.6000 12.2000 92.9000 13.8000 ;
	    RECT 93.4000 12.4000 93.8000 13.2000 ;
	    RECT 95.0000 12.2000 95.3000 13.8000 ;
	    RECT 95.8000 13.2000 96.1000 13.8000 ;
	    RECT 95.8000 13.1000 96.2000 13.2000 ;
	    RECT 97.4000 13.1000 97.8000 19.9000 ;
	    RECT 100.6000 16.2000 101.0000 19.9000 ;
	    RECT 102.2000 16.2000 102.6000 19.9000 ;
	    RECT 100.6000 15.9000 102.6000 16.2000 ;
	    RECT 103.0000 15.9000 103.4000 19.9000 ;
	    RECT 105.1000 16.3000 105.5000 19.9000 ;
	    RECT 107.5000 16.3000 107.9000 19.9000 ;
	    RECT 104.6000 15.9000 105.5000 16.3000 ;
	    RECT 107.0000 15.9000 107.9000 16.3000 ;
	    RECT 108.6000 15.9000 109.0000 19.9000 ;
	    RECT 109.4000 16.2000 109.8000 19.9000 ;
	    RECT 111.0000 16.2000 111.4000 19.9000 ;
	    RECT 112.6000 16.4000 113.0000 19.9000 ;
	    RECT 109.4000 15.9000 111.4000 16.2000 ;
	    RECT 112.5000 15.9000 113.0000 16.4000 ;
	    RECT 114.2000 16.2000 114.6000 19.9000 ;
	    RECT 113.3000 15.9000 114.6000 16.2000 ;
	    RECT 115.0000 16.2000 115.4000 19.9000 ;
	    RECT 116.6000 16.4000 117.0000 19.9000 ;
	    RECT 119.0000 16.4000 119.4000 19.9000 ;
	    RECT 115.0000 15.9000 116.3000 16.2000 ;
	    RECT 116.6000 15.9000 117.1000 16.4000 ;
	    RECT 101.0000 15.2000 101.4000 15.4000 ;
	    RECT 103.0000 15.2000 103.3000 15.9000 ;
	    RECT 100.6000 14.9000 101.4000 15.2000 ;
	    RECT 102.2000 14.9000 103.4000 15.2000 ;
	    RECT 100.6000 14.8000 101.0000 14.9000 ;
	    RECT 98.2000 13.4000 98.6000 14.2000 ;
	    RECT 101.4000 13.8000 101.8000 14.6000 ;
	    RECT 95.8000 12.8000 97.8000 13.1000 ;
	    RECT 102.2000 13.1000 102.5000 14.9000 ;
	    RECT 103.0000 14.8000 103.4000 14.9000 ;
	    RECT 104.7000 14.2000 105.0000 15.9000 ;
	    RECT 105.4000 14.8000 105.8000 15.6000 ;
	    RECT 107.1000 14.2000 107.4000 15.9000 ;
	    RECT 107.8000 14.8000 108.2000 15.6000 ;
	    RECT 108.7000 15.2000 109.0000 15.9000 ;
	    RECT 110.6000 15.2000 111.0000 15.4000 ;
	    RECT 108.6000 14.9000 109.8000 15.2000 ;
	    RECT 110.6000 14.9000 111.4000 15.2000 ;
	    RECT 108.6000 14.8000 109.0000 14.9000 ;
	    RECT 104.6000 14.1000 105.0000 14.2000 ;
	    RECT 103.0000 13.8000 105.0000 14.1000 ;
	    RECT 107.0000 13.8000 107.4000 14.2000 ;
	    RECT 108.6000 14.1000 109.0000 14.2000 ;
	    RECT 109.5000 14.1000 109.8000 14.9000 ;
	    RECT 111.0000 14.8000 111.4000 14.9000 ;
	    RECT 108.6000 13.8000 109.8000 14.1000 ;
	    RECT 110.2000 14.1000 110.6000 14.6000 ;
	    RECT 112.5000 14.2000 112.8000 15.9000 ;
	    RECT 113.3000 14.9000 113.6000 15.9000 ;
	    RECT 113.1000 14.5000 113.6000 14.9000 ;
	    RECT 112.5000 14.1000 113.0000 14.2000 ;
	    RECT 110.2000 13.8000 113.0000 14.1000 ;
	    RECT 103.0000 13.2000 103.3000 13.8000 ;
	    RECT 95.8000 12.4000 96.2000 12.8000 ;
	    RECT 87.0000 11.1000 87.4000 11.8000 ;
	    RECT 88.6000 11.1000 89.0000 12.1000 ;
	    RECT 92.6000 11.1000 93.0000 12.2000 ;
	    RECT 95.0000 11.1000 95.4000 12.2000 ;
	    RECT 96.9000 11.1000 97.3000 12.8000 ;
	    RECT 102.2000 11.1000 102.6000 13.1000 ;
	    RECT 103.0000 12.8000 103.4000 13.2000 ;
	    RECT 102.9000 12.4000 103.3000 12.8000 ;
	    RECT 103.8000 12.4000 104.2000 13.2000 ;
	    RECT 104.7000 12.1000 105.0000 13.8000 ;
	    RECT 106.2000 12.4000 106.6000 13.2000 ;
	    RECT 107.1000 13.1000 107.4000 13.8000 ;
	    RECT 108.6000 13.1000 109.0000 13.2000 ;
	    RECT 109.5000 13.1000 109.8000 13.8000 ;
	    RECT 107.0000 12.8000 109.0000 13.1000 ;
	    RECT 107.1000 12.1000 107.4000 12.8000 ;
	    RECT 108.7000 12.4000 109.1000 12.8000 ;
	    RECT 104.6000 11.1000 105.0000 12.1000 ;
	    RECT 107.0000 11.1000 107.4000 12.1000 ;
	    RECT 109.4000 11.1000 109.8000 13.1000 ;
	    RECT 112.5000 13.1000 112.8000 13.8000 ;
	    RECT 113.3000 13.7000 113.6000 14.5000 ;
	    RECT 114.1000 15.1000 114.6000 15.2000 ;
	    RECT 115.0000 15.1000 115.5000 15.2000 ;
	    RECT 114.1000 14.8000 115.5000 15.1000 ;
	    RECT 114.1000 14.4000 114.5000 14.8000 ;
	    RECT 115.1000 14.4000 115.5000 14.8000 ;
	    RECT 116.0000 14.9000 116.3000 15.9000 ;
	    RECT 116.0000 14.5000 116.5000 14.9000 ;
	    RECT 116.0000 13.7000 116.3000 14.5000 ;
	    RECT 116.8000 14.2000 117.1000 15.9000 ;
	    RECT 118.9000 15.9000 119.4000 16.4000 ;
	    RECT 120.6000 16.2000 121.0000 19.9000 ;
	    RECT 119.7000 15.9000 121.0000 16.2000 ;
	    RECT 121.7000 16.3000 122.1000 19.9000 ;
	    RECT 121.7000 15.9000 122.6000 16.3000 ;
	    RECT 118.9000 14.2000 119.2000 15.9000 ;
	    RECT 119.7000 14.9000 120.0000 15.9000 ;
	    RECT 119.5000 14.5000 120.0000 14.9000 ;
	    RECT 116.6000 14.1000 117.1000 14.2000 ;
	    RECT 117.4000 14.1000 117.8000 14.2000 ;
	    RECT 116.6000 13.8000 117.8000 14.1000 ;
	    RECT 118.9000 13.8000 119.4000 14.2000 ;
	    RECT 113.3000 13.4000 114.6000 13.7000 ;
	    RECT 112.5000 12.8000 113.0000 13.1000 ;
	    RECT 112.6000 11.1000 113.0000 12.8000 ;
	    RECT 114.2000 11.1000 114.6000 13.4000 ;
	    RECT 115.0000 13.4000 116.3000 13.7000 ;
	    RECT 115.0000 11.1000 115.4000 13.4000 ;
	    RECT 116.8000 13.1000 117.1000 13.8000 ;
	    RECT 116.6000 12.8000 117.1000 13.1000 ;
	    RECT 118.9000 13.1000 119.2000 13.8000 ;
	    RECT 119.7000 13.7000 120.0000 14.5000 ;
	    RECT 120.5000 14.8000 121.0000 15.2000 ;
	    RECT 121.4000 14.8000 121.8000 15.6000 ;
	    RECT 122.2000 15.1000 122.5000 15.9000 ;
	    RECT 122.2000 14.8000 123.3000 15.1000 ;
	    RECT 120.5000 14.4000 120.9000 14.8000 ;
	    RECT 122.2000 14.2000 122.5000 14.8000 ;
	    RECT 123.0000 14.2000 123.3000 14.8000 ;
	    RECT 122.2000 13.8000 122.6000 14.2000 ;
	    RECT 123.0000 13.8000 123.4000 14.2000 ;
	    RECT 119.7000 13.4000 121.0000 13.7000 ;
	    RECT 118.9000 12.8000 119.4000 13.1000 ;
	    RECT 116.6000 11.1000 117.0000 12.8000 ;
	    RECT 119.0000 11.1000 119.4000 12.8000 ;
	    RECT 120.6000 11.1000 121.0000 13.4000 ;
	    RECT 122.2000 12.1000 122.5000 13.8000 ;
	    RECT 123.0000 13.1000 123.4000 13.2000 ;
	    RECT 123.8000 13.1000 124.2000 19.9000 ;
	    RECT 124.6000 17.1000 125.0000 17.2000 ;
	    RECT 125.4000 17.1000 125.8000 19.9000 ;
	    RECT 127.5000 17.9000 128.1000 19.9000 ;
	    RECT 129.8000 17.9000 130.2000 19.9000 ;
	    RECT 132.0000 18.2000 132.4000 19.9000 ;
	    RECT 132.0000 17.9000 133.0000 18.2000 ;
	    RECT 127.8000 17.5000 128.2000 17.9000 ;
	    RECT 129.9000 17.6000 130.2000 17.9000 ;
	    RECT 129.5000 17.3000 131.3000 17.6000 ;
	    RECT 132.6000 17.5000 133.0000 17.9000 ;
	    RECT 129.5000 17.2000 129.9000 17.3000 ;
	    RECT 130.9000 17.2000 131.3000 17.3000 ;
	    RECT 124.6000 16.8000 125.8000 17.1000 ;
	    RECT 125.4000 15.6000 125.8000 16.8000 ;
	    RECT 127.4000 16.6000 128.1000 17.0000 ;
	    RECT 127.8000 16.1000 128.1000 16.6000 ;
	    RECT 128.9000 16.5000 130.0000 16.8000 ;
	    RECT 128.9000 16.4000 129.3000 16.5000 ;
	    RECT 127.8000 15.8000 129.0000 16.1000 ;
	    RECT 125.4000 15.3000 127.5000 15.6000 ;
	    RECT 125.4000 13.6000 125.8000 15.3000 ;
	    RECT 127.1000 15.2000 127.5000 15.3000 ;
	    RECT 126.3000 14.9000 126.7000 15.0000 ;
	    RECT 126.3000 14.6000 128.2000 14.9000 ;
	    RECT 127.8000 14.5000 128.2000 14.6000 ;
	    RECT 128.7000 14.2000 129.0000 15.8000 ;
	    RECT 129.7000 15.9000 130.0000 16.5000 ;
	    RECT 130.3000 16.5000 130.7000 16.6000 ;
	    RECT 132.6000 16.5000 133.0000 16.6000 ;
	    RECT 130.3000 16.2000 133.0000 16.5000 ;
	    RECT 129.7000 15.7000 132.1000 15.9000 ;
	    RECT 134.2000 15.7000 134.6000 19.9000 ;
	    RECT 129.7000 15.6000 134.6000 15.7000 ;
	    RECT 131.7000 15.5000 134.6000 15.6000 ;
	    RECT 131.8000 15.4000 134.6000 15.5000 ;
	    RECT 135.0000 15.7000 135.4000 19.9000 ;
	    RECT 137.2000 18.2000 137.6000 19.9000 ;
	    RECT 136.6000 17.9000 137.6000 18.2000 ;
	    RECT 139.4000 17.9000 139.8000 19.9000 ;
	    RECT 141.5000 17.9000 142.1000 19.9000 ;
	    RECT 136.6000 17.5000 137.0000 17.9000 ;
	    RECT 139.4000 17.6000 139.7000 17.9000 ;
	    RECT 138.3000 17.3000 140.1000 17.6000 ;
	    RECT 141.4000 17.5000 141.8000 17.9000 ;
	    RECT 138.3000 17.2000 138.7000 17.3000 ;
	    RECT 139.7000 17.2000 140.1000 17.3000 ;
	    RECT 136.6000 16.5000 137.0000 16.6000 ;
	    RECT 138.9000 16.5000 139.3000 16.6000 ;
	    RECT 136.6000 16.2000 139.3000 16.5000 ;
	    RECT 139.6000 16.5000 140.7000 16.8000 ;
	    RECT 139.6000 15.9000 139.9000 16.5000 ;
	    RECT 140.3000 16.4000 140.7000 16.5000 ;
	    RECT 141.5000 16.6000 142.2000 17.0000 ;
	    RECT 141.5000 16.1000 141.8000 16.6000 ;
	    RECT 137.5000 15.7000 139.9000 15.9000 ;
	    RECT 135.0000 15.6000 139.9000 15.7000 ;
	    RECT 140.6000 15.8000 141.8000 16.1000 ;
	    RECT 135.0000 15.5000 137.9000 15.6000 ;
	    RECT 135.0000 15.4000 137.8000 15.5000 ;
	    RECT 129.4000 15.1000 129.8000 15.2000 ;
	    RECT 131.0000 15.1000 131.4000 15.2000 ;
	    RECT 138.2000 15.1000 138.6000 15.2000 ;
	    RECT 129.4000 14.8000 133.5000 15.1000 ;
	    RECT 133.1000 14.7000 133.5000 14.8000 ;
	    RECT 136.1000 14.8000 138.6000 15.1000 ;
	    RECT 136.1000 14.7000 136.5000 14.8000 ;
	    RECT 137.4000 14.7000 137.8000 14.8000 ;
	    RECT 132.3000 14.2000 132.7000 14.3000 ;
	    RECT 136.9000 14.2000 137.3000 14.3000 ;
	    RECT 140.6000 14.2000 140.9000 15.8000 ;
	    RECT 143.8000 15.6000 144.2000 19.9000 ;
	    RECT 144.6000 16.2000 145.0000 19.9000 ;
	    RECT 146.2000 16.4000 146.6000 19.9000 ;
	    RECT 144.6000 15.9000 145.9000 16.2000 ;
	    RECT 146.2000 15.9000 146.7000 16.4000 ;
	    RECT 142.1000 15.3000 144.2000 15.6000 ;
	    RECT 142.1000 15.2000 142.5000 15.3000 ;
	    RECT 142.9000 14.9000 143.3000 15.0000 ;
	    RECT 141.4000 14.6000 143.3000 14.9000 ;
	    RECT 141.4000 14.5000 141.8000 14.6000 ;
	    RECT 128.7000 14.1000 134.2000 14.2000 ;
	    RECT 135.4000 14.1000 140.9000 14.2000 ;
	    RECT 128.7000 13.9000 140.9000 14.1000 ;
	    RECT 128.9000 13.8000 129.3000 13.9000 ;
	    RECT 125.4000 13.3000 127.3000 13.6000 ;
	    RECT 123.0000 12.8000 124.2000 13.1000 ;
	    RECT 123.0000 12.4000 123.4000 12.8000 ;
	    RECT 122.2000 11.1000 122.6000 12.1000 ;
	    RECT 123.8000 11.1000 124.2000 12.8000 ;
	    RECT 124.6000 12.4000 125.0000 13.2000 ;
	    RECT 125.4000 11.1000 125.8000 13.3000 ;
	    RECT 126.9000 13.2000 127.3000 13.3000 ;
	    RECT 131.8000 12.8000 132.1000 13.9000 ;
	    RECT 133.4000 13.8000 136.2000 13.9000 ;
	    RECT 130.9000 12.7000 131.3000 12.8000 ;
	    RECT 127.8000 12.1000 128.2000 12.5000 ;
	    RECT 129.9000 12.4000 131.3000 12.7000 ;
	    RECT 131.8000 12.4000 132.2000 12.8000 ;
	    RECT 129.9000 12.1000 130.2000 12.4000 ;
	    RECT 132.6000 12.1000 133.0000 12.5000 ;
	    RECT 127.5000 11.8000 128.2000 12.1000 ;
	    RECT 127.5000 11.1000 128.1000 11.8000 ;
	    RECT 129.8000 11.1000 130.2000 12.1000 ;
	    RECT 132.0000 11.8000 133.0000 12.1000 ;
	    RECT 132.0000 11.1000 132.4000 11.8000 ;
	    RECT 134.2000 11.1000 134.6000 13.5000 ;
	    RECT 135.0000 11.1000 135.4000 13.5000 ;
	    RECT 137.5000 12.8000 137.8000 13.9000 ;
	    RECT 138.2000 13.8000 138.6000 13.9000 ;
	    RECT 140.3000 13.8000 140.7000 13.9000 ;
	    RECT 143.8000 13.6000 144.2000 15.3000 ;
	    RECT 144.6000 14.8000 145.1000 15.2000 ;
	    RECT 144.7000 14.4000 145.1000 14.8000 ;
	    RECT 145.6000 14.9000 145.9000 15.9000 ;
	    RECT 145.6000 14.5000 146.1000 14.9000 ;
	    RECT 145.6000 13.7000 145.9000 14.5000 ;
	    RECT 146.4000 14.2000 146.7000 15.9000 ;
	    RECT 146.2000 13.8000 146.7000 14.2000 ;
	    RECT 142.3000 13.3000 144.2000 13.6000 ;
	    RECT 142.3000 13.2000 142.7000 13.3000 ;
	    RECT 136.6000 12.1000 137.0000 12.5000 ;
	    RECT 137.4000 12.4000 137.8000 12.8000 ;
	    RECT 138.3000 12.7000 138.7000 12.8000 ;
	    RECT 138.3000 12.4000 139.7000 12.7000 ;
	    RECT 139.4000 12.1000 139.7000 12.4000 ;
	    RECT 141.4000 12.1000 141.8000 12.5000 ;
	    RECT 136.6000 11.8000 137.6000 12.1000 ;
	    RECT 137.2000 11.1000 137.6000 11.8000 ;
	    RECT 139.4000 11.1000 139.8000 12.1000 ;
	    RECT 141.4000 11.8000 142.1000 12.1000 ;
	    RECT 141.5000 11.1000 142.1000 11.8000 ;
	    RECT 143.8000 11.1000 144.2000 13.3000 ;
	    RECT 144.6000 13.4000 145.9000 13.7000 ;
	    RECT 144.6000 11.1000 145.0000 13.4000 ;
	    RECT 146.4000 13.1000 146.7000 13.8000 ;
	    RECT 146.2000 12.8000 146.7000 13.1000 ;
	    RECT 146.2000 11.1000 146.6000 12.8000 ;
	    RECT 2.2000 7.6000 2.6000 9.9000 ;
	    RECT 1.5000 7.3000 2.6000 7.6000 ;
	    RECT 1.5000 5.8000 1.8000 7.3000 ;
	    RECT 3.8000 7.1000 4.2000 9.9000 ;
	    RECT 6.2000 7.9000 6.6000 9.9000 ;
	    RECT 8.6000 8.9000 9.0000 9.9000 ;
	    RECT 6.9000 8.2000 7.3000 8.6000 ;
	    RECT 4.6000 7.1000 5.0000 7.2000 ;
	    RECT 3.8000 6.8000 5.0000 7.1000 ;
	    RECT 2.2000 5.8000 2.6000 6.6000 ;
	    RECT 3.8000 6.1000 4.2000 6.8000 ;
	    RECT 5.4000 6.4000 5.8000 7.2000 ;
	    RECT 4.6000 6.1000 5.0000 6.2000 ;
	    RECT 6.2000 6.1000 6.5000 7.9000 ;
	    RECT 7.0000 7.8000 7.4000 8.2000 ;
	    RECT 7.8000 7.8000 8.2000 8.6000 ;
	    RECT 8.7000 7.2000 9.0000 8.9000 ;
	    RECT 10.5000 8.2000 10.9000 9.9000 ;
	    RECT 15.0000 8.9000 15.4000 9.9000 ;
	    RECT 16.6000 9.2000 17.0000 9.9000 ;
	    RECT 14.8000 8.8000 15.4000 8.9000 ;
	    RECT 16.5000 8.8000 17.0000 9.2000 ;
	    RECT 19.8000 8.9000 20.2000 9.9000 ;
	    RECT 23.0000 9.2000 23.4000 9.9000 ;
	    RECT 23.0000 8.9000 23.5000 9.2000 ;
	    RECT 14.8000 8.5000 16.8000 8.8000 ;
	    RECT 7.8000 6.8000 8.2000 7.2000 ;
	    RECT 8.6000 6.8000 9.0000 7.2000 ;
	    RECT 10.2000 7.8000 11.4000 8.2000 ;
	    RECT 10.2000 7.2000 10.5000 7.8000 ;
	    RECT 10.2000 6.8000 10.6000 7.2000 ;
	    RECT 7.0000 6.1000 7.4000 6.2000 ;
	    RECT 3.8000 5.8000 5.4000 6.1000 ;
	    RECT 6.2000 5.8000 7.4000 6.1000 ;
	    RECT 7.8000 6.1000 8.1000 6.8000 ;
	    RECT 8.7000 6.1000 9.0000 6.8000 ;
	    RECT 7.8000 5.8000 9.0000 6.1000 ;
	    RECT 1.2000 5.4000 1.8000 5.8000 ;
	    RECT 1.5000 5.1000 1.8000 5.4000 ;
	    RECT 1.5000 4.8000 2.6000 5.1000 ;
	    RECT 2.2000 1.1000 2.6000 4.8000 ;
	    RECT 3.8000 1.1000 4.2000 5.8000 ;
	    RECT 5.0000 5.6000 5.4000 5.8000 ;
	    RECT 7.0000 5.1000 7.3000 5.8000 ;
	    RECT 8.7000 5.1000 9.0000 5.8000 ;
	    RECT 9.4000 5.4000 9.8000 6.2000 ;
	    RECT 4.6000 4.8000 6.6000 5.1000 ;
	    RECT 4.6000 1.1000 5.0000 4.8000 ;
	    RECT 6.2000 1.1000 6.6000 4.8000 ;
	    RECT 7.0000 1.1000 7.4000 5.1000 ;
	    RECT 8.6000 4.7000 9.5000 5.1000 ;
	    RECT 9.1000 1.1000 9.5000 4.7000 ;
	    RECT 10.2000 4.4000 10.6000 5.2000 ;
	    RECT 11.0000 1.1000 11.4000 7.8000 ;
	    RECT 11.8000 6.8000 12.2000 7.6000 ;
	    RECT 14.8000 5.2000 15.1000 8.5000 ;
	    RECT 16.6000 7.8000 17.8000 8.2000 ;
	    RECT 19.8000 7.2000 20.1000 8.9000 ;
	    RECT 23.2000 8.8000 23.5000 8.9000 ;
	    RECT 24.6000 9.1000 25.0000 9.9000 ;
	    RECT 27.0000 9.1000 27.4000 9.2000 ;
	    RECT 24.6000 8.8000 27.4000 9.1000 ;
	    RECT 23.2000 8.5000 25.2000 8.8000 ;
	    RECT 22.2000 7.8000 23.1000 8.2000 ;
	    RECT 16.2000 7.1000 17.0000 7.2000 ;
	    RECT 18.2000 7.1000 18.6000 7.2000 ;
	    RECT 16.2000 6.8000 18.6000 7.1000 ;
	    RECT 19.8000 6.8000 20.2000 7.2000 ;
	    RECT 23.0000 6.8000 23.8000 7.2000 ;
	    RECT 15.4000 5.8000 16.2000 6.2000 ;
	    RECT 19.0000 5.4000 19.4000 6.2000 ;
	    RECT 13.4000 4.9000 15.1000 5.2000 ;
	    RECT 19.8000 5.1000 20.1000 6.8000 ;
	    RECT 23.8000 5.8000 24.6000 6.2000 ;
	    RECT 24.9000 5.2000 25.2000 8.5000 ;
	    RECT 27.8000 6.8000 28.2000 7.6000 ;
	    RECT 28.6000 6.1000 29.0000 9.9000 ;
	    RECT 29.4000 8.0000 29.8000 9.9000 ;
	    RECT 31.0000 8.0000 31.4000 9.9000 ;
	    RECT 29.4000 7.9000 31.4000 8.0000 ;
	    RECT 31.8000 7.9000 32.2000 9.9000 ;
	    RECT 32.6000 7.9000 33.0000 9.9000 ;
	    RECT 33.4000 8.0000 33.8000 9.9000 ;
	    RECT 35.0000 8.0000 35.4000 9.9000 ;
	    RECT 37.4000 9.2000 37.8000 9.9000 ;
	    RECT 37.4000 8.8000 37.9000 9.2000 ;
	    RECT 39.0000 8.9000 39.4000 9.9000 ;
	    RECT 43.0000 9.1000 43.4000 9.2000 ;
	    RECT 44.0000 9.1000 44.4000 9.9000 ;
	    RECT 39.0000 8.8000 39.6000 8.9000 ;
	    RECT 43.0000 8.8000 44.4000 9.1000 ;
	    RECT 37.6000 8.5000 39.6000 8.8000 ;
	    RECT 33.4000 7.9000 35.4000 8.0000 ;
	    RECT 29.5000 7.7000 31.3000 7.9000 ;
	    RECT 29.8000 7.2000 30.2000 7.4000 ;
	    RECT 31.8000 7.2000 32.1000 7.9000 ;
	    RECT 32.7000 7.2000 33.0000 7.9000 ;
	    RECT 33.5000 7.7000 35.3000 7.9000 ;
	    RECT 34.6000 7.2000 35.0000 7.4000 ;
	    RECT 29.4000 6.9000 30.2000 7.2000 ;
	    RECT 29.4000 6.8000 29.8000 6.9000 ;
	    RECT 30.9000 6.8000 32.2000 7.2000 ;
	    RECT 32.6000 6.8000 33.9000 7.2000 ;
	    RECT 34.6000 6.9000 35.4000 7.2000 ;
	    RECT 37.4000 7.1000 38.2000 7.2000 ;
	    RECT 35.0000 6.8000 35.4000 6.9000 ;
	    RECT 35.8000 6.8000 38.2000 7.1000 ;
	    RECT 30.2000 6.1000 30.6000 6.6000 ;
	    RECT 28.6000 5.8000 30.6000 6.1000 ;
	    RECT 13.4000 4.8000 13.8000 4.9000 ;
	    RECT 13.5000 4.5000 13.8000 4.8000 ;
	    RECT 19.3000 4.7000 20.2000 5.1000 ;
	    RECT 24.9000 4.9000 26.6000 5.2000 ;
	    RECT 26.2000 4.8000 26.6000 4.9000 ;
	    RECT 14.3000 4.5000 16.1000 4.6000 ;
	    RECT 12.6000 1.5000 13.0000 4.5000 ;
	    RECT 13.4000 1.7000 13.8000 4.5000 ;
	    RECT 14.2000 4.3000 16.1000 4.5000 ;
	    RECT 12.7000 1.4000 13.0000 1.5000 ;
	    RECT 14.2000 1.5000 14.6000 4.3000 ;
	    RECT 15.8000 4.1000 16.1000 4.3000 ;
	    RECT 16.7000 4.4000 18.5000 4.7000 ;
	    RECT 16.7000 4.1000 17.0000 4.4000 ;
	    RECT 14.2000 1.4000 14.5000 1.5000 ;
	    RECT 12.7000 1.1000 14.5000 1.4000 ;
	    RECT 15.0000 1.4000 15.4000 4.0000 ;
	    RECT 15.8000 1.7000 16.2000 4.1000 ;
	    RECT 16.6000 1.4000 17.0000 4.1000 ;
	    RECT 15.0000 1.1000 17.0000 1.4000 ;
	    RECT 18.2000 4.1000 18.5000 4.4000 ;
	    RECT 19.3000 4.2000 19.7000 4.7000 ;
	    RECT 18.2000 1.1000 18.6000 4.1000 ;
	    RECT 19.0000 3.8000 19.7000 4.2000 ;
	    RECT 21.5000 4.4000 23.3000 4.7000 ;
	    RECT 21.5000 4.1000 21.8000 4.4000 ;
	    RECT 19.3000 1.1000 19.7000 3.8000 ;
	    RECT 21.4000 1.1000 21.8000 4.1000 ;
	    RECT 23.0000 4.1000 23.3000 4.4000 ;
	    RECT 23.9000 4.5000 25.7000 4.6000 ;
	    RECT 26.2000 4.5000 26.5000 4.8000 ;
	    RECT 23.9000 4.3000 25.8000 4.5000 ;
	    RECT 23.9000 4.1000 24.2000 4.3000 ;
	    RECT 23.0000 1.4000 23.4000 4.1000 ;
	    RECT 23.8000 1.7000 24.2000 4.1000 ;
	    RECT 24.6000 1.4000 25.0000 4.0000 ;
	    RECT 25.4000 1.5000 25.8000 4.3000 ;
	    RECT 26.2000 1.7000 26.6000 4.5000 ;
	    RECT 23.0000 1.1000 25.0000 1.4000 ;
	    RECT 25.5000 1.4000 25.8000 1.5000 ;
	    RECT 27.0000 1.5000 27.4000 4.5000 ;
	    RECT 27.0000 1.4000 27.3000 1.5000 ;
	    RECT 25.5000 1.1000 27.3000 1.4000 ;
	    RECT 28.6000 1.1000 29.0000 5.8000 ;
	    RECT 30.9000 5.2000 31.2000 6.8000 ;
	    RECT 33.6000 6.1000 33.9000 6.8000 ;
	    RECT 30.8000 5.1000 31.2000 5.2000 ;
	    RECT 31.8000 5.8000 33.9000 6.1000 ;
	    RECT 34.2000 6.1000 34.6000 6.6000 ;
	    RECT 35.8000 6.1000 36.1000 6.8000 ;
	    RECT 34.2000 5.8000 36.1000 6.1000 ;
	    RECT 38.2000 5.8000 39.0000 6.2000 ;
	    RECT 31.8000 5.2000 32.1000 5.8000 ;
	    RECT 31.8000 5.1000 32.2000 5.2000 ;
	    RECT 30.7000 4.8000 31.2000 5.1000 ;
	    RECT 31.5000 4.8000 32.2000 5.1000 ;
	    RECT 32.6000 5.1000 33.0000 5.2000 ;
	    RECT 33.6000 5.1000 33.9000 5.8000 ;
	    RECT 39.3000 5.2000 39.6000 8.5000 ;
	    RECT 44.0000 7.1000 44.4000 8.8000 ;
	    RECT 46.2000 8.9000 46.6000 9.9000 ;
	    RECT 46.2000 7.2000 46.5000 8.9000 ;
	    RECT 47.0000 7.8000 47.4000 8.6000 ;
	    RECT 49.4000 8.0000 49.8000 9.9000 ;
	    RECT 51.0000 8.0000 51.4000 9.9000 ;
	    RECT 49.4000 7.9000 51.4000 8.0000 ;
	    RECT 51.8000 7.9000 52.2000 9.9000 ;
	    RECT 54.2000 9.2000 54.6000 9.9000 ;
	    RECT 54.2000 8.9000 54.7000 9.2000 ;
	    RECT 54.4000 8.8000 54.7000 8.9000 ;
	    RECT 55.8000 8.9000 56.2000 9.9000 ;
	    RECT 55.8000 8.8000 56.4000 8.9000 ;
	    RECT 54.4000 8.5000 56.4000 8.8000 ;
	    RECT 49.5000 7.7000 51.3000 7.9000 ;
	    RECT 49.8000 7.2000 50.2000 7.4000 ;
	    RECT 51.8000 7.2000 52.1000 7.9000 ;
	    RECT 53.4000 7.8000 54.3000 8.2000 ;
	    RECT 44.0000 6.9000 44.9000 7.1000 ;
	    RECT 44.1000 6.8000 44.9000 6.9000 ;
	    RECT 43.0000 5.8000 43.8000 6.2000 ;
	    RECT 44.6000 6.1000 44.9000 6.8000 ;
	    RECT 46.2000 6.8000 46.6000 7.2000 ;
	    RECT 49.4000 6.9000 50.2000 7.2000 ;
	    RECT 49.4000 6.8000 49.8000 6.9000 ;
	    RECT 50.9000 6.8000 52.2000 7.2000 ;
	    RECT 53.4000 7.1000 53.8000 7.2000 ;
	    RECT 54.2000 7.1000 55.0000 7.2000 ;
	    RECT 53.4000 6.8000 55.0000 7.1000 ;
	    RECT 46.2000 6.2000 46.5000 6.8000 ;
	    RECT 45.4000 6.1000 45.8000 6.2000 ;
	    RECT 44.6000 5.8000 45.8000 6.1000 ;
	    RECT 44.6000 5.2000 44.9000 5.8000 ;
	    RECT 45.4000 5.4000 45.8000 5.8000 ;
	    RECT 46.2000 5.8000 46.6000 6.2000 ;
	    RECT 47.0000 6.1000 47.4000 6.2000 ;
	    RECT 50.2000 6.1000 50.6000 6.6000 ;
	    RECT 47.0000 5.8000 50.6000 6.1000 ;
	    RECT 32.6000 4.8000 33.3000 5.1000 ;
	    RECT 33.6000 4.8000 34.1000 5.1000 ;
	    RECT 39.3000 4.9000 41.0000 5.2000 ;
	    RECT 30.7000 1.1000 31.1000 4.8000 ;
	    RECT 31.5000 4.2000 31.8000 4.8000 ;
	    RECT 31.4000 3.8000 31.8000 4.2000 ;
	    RECT 33.0000 4.2000 33.3000 4.8000 ;
	    RECT 33.0000 3.8000 33.4000 4.2000 ;
	    RECT 33.7000 1.1000 34.1000 4.8000 ;
	    RECT 40.6000 4.8000 41.0000 4.9000 ;
	    RECT 44.6000 4.8000 45.0000 5.2000 ;
	    RECT 46.2000 5.1000 46.5000 5.8000 ;
	    RECT 50.9000 5.2000 51.2000 6.8000 ;
	    RECT 52.6000 6.1000 53.0000 6.2000 ;
	    RECT 50.8000 5.1000 51.2000 5.2000 ;
	    RECT 51.8000 5.8000 53.0000 6.1000 ;
	    RECT 55.0000 5.8000 55.8000 6.2000 ;
	    RECT 51.8000 5.2000 52.1000 5.8000 ;
	    RECT 56.1000 5.2000 56.4000 8.5000 ;
	    RECT 59.0000 8.0000 59.4000 9.9000 ;
	    RECT 60.6000 8.0000 61.0000 9.9000 ;
	    RECT 59.0000 7.9000 61.0000 8.0000 ;
	    RECT 61.4000 7.9000 61.8000 9.9000 ;
	    RECT 62.5000 8.2000 62.9000 9.9000 ;
	    RECT 62.5000 7.9000 63.4000 8.2000 ;
	    RECT 59.1000 7.7000 60.9000 7.9000 ;
	    RECT 59.4000 7.2000 59.8000 7.4000 ;
	    RECT 61.4000 7.2000 61.7000 7.9000 ;
	    RECT 59.0000 6.9000 59.8000 7.2000 ;
	    RECT 59.0000 6.8000 59.4000 6.9000 ;
	    RECT 60.5000 6.8000 61.8000 7.2000 ;
	    RECT 62.2000 6.8000 62.6000 7.2000 ;
	    RECT 58.2000 6.1000 58.6000 6.2000 ;
	    RECT 59.8000 6.1000 60.2000 6.6000 ;
	    RECT 58.2000 5.8000 60.2000 6.1000 ;
	    RECT 60.5000 6.1000 60.8000 6.8000 ;
	    RECT 62.2000 6.1000 62.5000 6.8000 ;
	    RECT 60.5000 5.8000 62.5000 6.1000 ;
	    RECT 51.8000 5.1000 52.2000 5.2000 ;
	    RECT 35.9000 4.4000 37.7000 4.7000 ;
	    RECT 35.9000 4.1000 36.2000 4.4000 ;
	    RECT 35.8000 1.1000 36.2000 4.1000 ;
	    RECT 37.4000 4.1000 37.7000 4.4000 ;
	    RECT 38.3000 4.5000 40.1000 4.6000 ;
	    RECT 40.6000 4.5000 40.9000 4.8000 ;
	    RECT 38.3000 4.3000 40.2000 4.5000 ;
	    RECT 38.3000 4.1000 38.6000 4.3000 ;
	    RECT 37.4000 1.4000 37.8000 4.1000 ;
	    RECT 38.2000 1.7000 38.6000 4.1000 ;
	    RECT 39.0000 1.4000 39.4000 4.0000 ;
	    RECT 39.8000 1.5000 40.2000 4.3000 ;
	    RECT 40.6000 1.7000 41.0000 4.5000 ;
	    RECT 37.4000 1.1000 39.4000 1.4000 ;
	    RECT 39.9000 1.4000 40.2000 1.5000 ;
	    RECT 41.4000 1.5000 41.8000 4.5000 ;
	    RECT 43.8000 3.8000 44.2000 4.6000 ;
	    RECT 44.6000 3.5000 44.9000 4.8000 ;
	    RECT 43.1000 3.2000 44.9000 3.5000 ;
	    RECT 43.1000 3.1000 43.4000 3.2000 ;
	    RECT 41.4000 1.4000 41.7000 1.5000 ;
	    RECT 39.9000 1.1000 41.7000 1.4000 ;
	    RECT 43.0000 1.1000 43.4000 3.1000 ;
	    RECT 44.6000 3.1000 44.9000 3.2000 ;
	    RECT 45.7000 4.7000 46.6000 5.1000 ;
	    RECT 50.7000 4.8000 51.2000 5.1000 ;
	    RECT 51.5000 4.8000 52.2000 5.1000 ;
	    RECT 56.1000 4.9000 57.8000 5.2000 ;
	    RECT 60.5000 5.1000 60.8000 5.8000 ;
	    RECT 57.4000 4.8000 57.8000 4.9000 ;
	    RECT 60.3000 4.8000 60.8000 5.1000 ;
	    RECT 44.6000 1.1000 45.0000 3.1000 ;
	    RECT 45.7000 1.1000 46.1000 4.7000 ;
	    RECT 50.7000 1.1000 51.1000 4.8000 ;
	    RECT 51.5000 4.2000 51.8000 4.8000 ;
	    RECT 51.4000 3.8000 51.8000 4.2000 ;
	    RECT 52.7000 4.4000 54.5000 4.7000 ;
	    RECT 52.7000 4.1000 53.0000 4.4000 ;
	    RECT 52.6000 1.1000 53.0000 4.1000 ;
	    RECT 54.2000 4.1000 54.5000 4.4000 ;
	    RECT 55.1000 4.5000 56.9000 4.6000 ;
	    RECT 57.4000 4.5000 57.7000 4.8000 ;
	    RECT 55.1000 4.3000 57.0000 4.5000 ;
	    RECT 55.1000 4.1000 55.4000 4.3000 ;
	    RECT 54.2000 1.4000 54.6000 4.1000 ;
	    RECT 55.0000 1.7000 55.4000 4.1000 ;
	    RECT 55.8000 1.4000 56.2000 4.0000 ;
	    RECT 56.6000 1.5000 57.0000 4.3000 ;
	    RECT 57.4000 1.7000 57.8000 4.5000 ;
	    RECT 54.2000 1.1000 56.2000 1.4000 ;
	    RECT 56.7000 1.4000 57.0000 1.5000 ;
	    RECT 58.2000 1.5000 58.6000 4.5000 ;
	    RECT 58.2000 1.4000 58.5000 1.5000 ;
	    RECT 56.7000 1.1000 58.5000 1.4000 ;
	    RECT 60.3000 1.1000 60.7000 4.8000 ;
	    RECT 62.2000 4.4000 62.6000 5.2000 ;
	    RECT 63.0000 5.1000 63.4000 7.9000 ;
	    RECT 64.6000 7.6000 65.0000 9.9000 ;
	    RECT 63.8000 6.8000 64.2000 7.6000 ;
	    RECT 64.6000 7.3000 65.7000 7.6000 ;
	    RECT 63.8000 5.8000 64.2000 6.2000 ;
	    RECT 64.6000 5.8000 65.0000 6.6000 ;
	    RECT 65.4000 5.8000 65.7000 7.3000 ;
	    RECT 68.8000 7.1000 69.2000 9.9000 ;
	    RECT 70.2000 7.7000 70.6000 9.9000 ;
	    RECT 72.3000 9.2000 72.9000 9.9000 ;
	    RECT 72.3000 8.9000 73.0000 9.2000 ;
	    RECT 74.6000 8.9000 75.0000 9.9000 ;
	    RECT 76.8000 9.2000 77.2000 9.9000 ;
	    RECT 76.8000 8.9000 77.8000 9.2000 ;
	    RECT 72.6000 8.5000 73.0000 8.9000 ;
	    RECT 74.7000 8.6000 75.0000 8.9000 ;
	    RECT 74.7000 8.3000 76.1000 8.6000 ;
	    RECT 75.7000 8.2000 76.1000 8.3000 ;
	    RECT 76.6000 8.2000 77.0000 8.6000 ;
	    RECT 77.4000 8.5000 77.8000 8.9000 ;
	    RECT 71.7000 7.7000 72.1000 7.8000 ;
	    RECT 70.2000 7.4000 72.1000 7.7000 ;
	    RECT 68.8000 6.9000 69.7000 7.1000 ;
	    RECT 68.9000 6.8000 69.7000 6.9000 ;
	    RECT 69.4000 6.2000 69.7000 6.8000 ;
	    RECT 67.8000 5.8000 68.6000 6.2000 ;
	    RECT 69.4000 5.8000 69.8000 6.2000 ;
	    RECT 63.8000 5.1000 64.1000 5.8000 ;
	    RECT 65.4000 5.4000 66.0000 5.8000 ;
	    RECT 65.4000 5.1000 65.7000 5.4000 ;
	    RECT 63.0000 4.8000 64.1000 5.1000 ;
	    RECT 64.6000 4.8000 65.7000 5.1000 ;
	    RECT 67.0000 4.8000 67.4000 5.6000 ;
	    RECT 69.4000 5.2000 69.7000 5.8000 ;
	    RECT 70.2000 5.7000 70.6000 7.4000 ;
	    RECT 73.7000 7.1000 74.1000 7.2000 ;
	    RECT 76.6000 7.1000 76.9000 8.2000 ;
	    RECT 79.0000 7.5000 79.4000 9.9000 ;
	    RECT 81.4000 7.6000 81.8000 9.9000 ;
	    RECT 83.8000 7.6000 84.2000 9.9000 ;
	    RECT 80.7000 7.3000 81.8000 7.6000 ;
	    RECT 83.1000 7.3000 84.2000 7.6000 ;
	    RECT 84.6000 7.5000 85.0000 9.9000 ;
	    RECT 86.8000 9.2000 87.2000 9.9000 ;
	    RECT 86.2000 8.9000 87.2000 9.2000 ;
	    RECT 89.0000 8.9000 89.4000 9.9000 ;
	    RECT 91.1000 9.2000 91.7000 9.9000 ;
	    RECT 91.0000 8.9000 91.7000 9.2000 ;
	    RECT 86.2000 8.5000 86.6000 8.9000 ;
	    RECT 89.0000 8.6000 89.3000 8.9000 ;
	    RECT 87.0000 8.2000 87.4000 8.6000 ;
	    RECT 87.9000 8.3000 89.3000 8.6000 ;
	    RECT 91.0000 8.5000 91.4000 8.9000 ;
	    RECT 87.9000 8.2000 88.3000 8.3000 ;
	    RECT 78.2000 7.1000 79.0000 7.2000 ;
	    RECT 73.5000 6.8000 79.0000 7.1000 ;
	    RECT 72.6000 6.4000 73.0000 6.5000 ;
	    RECT 71.1000 6.1000 73.0000 6.4000 ;
	    RECT 71.1000 6.0000 71.5000 6.1000 ;
	    RECT 71.9000 5.7000 72.3000 5.8000 ;
	    RECT 70.2000 5.4000 72.3000 5.7000 ;
	    RECT 69.4000 4.8000 69.8000 5.2000 ;
	    RECT 63.0000 1.1000 63.4000 4.8000 ;
	    RECT 64.6000 1.1000 65.0000 4.8000 ;
	    RECT 68.6000 3.8000 69.0000 4.6000 ;
	    RECT 69.4000 3.5000 69.7000 4.8000 ;
	    RECT 67.9000 3.2000 69.7000 3.5000 ;
	    RECT 67.9000 3.1000 68.2000 3.2000 ;
	    RECT 67.8000 1.1000 68.2000 3.1000 ;
	    RECT 69.4000 3.1000 69.7000 3.2000 ;
	    RECT 69.4000 1.1000 69.8000 3.1000 ;
	    RECT 70.2000 1.1000 70.6000 5.4000 ;
	    RECT 73.5000 5.2000 73.8000 6.8000 ;
	    RECT 77.1000 6.7000 77.5000 6.8000 ;
	    RECT 77.9000 6.2000 78.3000 6.3000 ;
	    RECT 75.8000 5.9000 78.3000 6.2000 ;
	    RECT 75.8000 5.8000 76.2000 5.9000 ;
	    RECT 80.7000 5.8000 81.0000 7.3000 ;
	    RECT 81.4000 5.8000 81.8000 6.6000 ;
	    RECT 83.1000 5.8000 83.4000 7.3000 ;
	    RECT 85.0000 7.1000 85.8000 7.2000 ;
	    RECT 87.1000 7.1000 87.4000 8.2000 ;
	    RECT 91.9000 7.7000 92.3000 7.8000 ;
	    RECT 93.4000 7.7000 93.8000 9.9000 ;
	    RECT 91.9000 7.4000 93.8000 7.7000 ;
	    RECT 89.9000 7.1000 90.3000 7.2000 ;
	    RECT 85.0000 6.8000 90.5000 7.1000 ;
	    RECT 86.5000 6.7000 86.9000 6.8000 ;
	    RECT 83.8000 5.8000 84.2000 6.6000 ;
	    RECT 85.7000 6.2000 86.1000 6.3000 ;
	    RECT 90.2000 6.2000 90.5000 6.8000 ;
	    RECT 91.0000 6.4000 91.4000 6.5000 ;
	    RECT 85.7000 5.9000 88.2000 6.2000 ;
	    RECT 87.8000 5.8000 88.2000 5.9000 ;
	    RECT 90.2000 5.8000 90.6000 6.2000 ;
	    RECT 91.0000 6.1000 92.9000 6.4000 ;
	    RECT 92.5000 6.0000 92.9000 6.1000 ;
	    RECT 93.4000 6.1000 93.8000 7.4000 ;
	    RECT 94.2000 7.6000 94.6000 9.9000 ;
	    RECT 96.6000 7.6000 97.0000 9.9000 ;
	    RECT 100.6000 7.7000 101.0000 9.9000 ;
	    RECT 102.7000 9.2000 103.3000 9.9000 ;
	    RECT 102.7000 8.9000 103.4000 9.2000 ;
	    RECT 105.0000 8.9000 105.4000 9.9000 ;
	    RECT 107.2000 9.2000 107.6000 9.9000 ;
	    RECT 107.2000 8.9000 108.2000 9.2000 ;
	    RECT 103.0000 8.5000 103.4000 8.9000 ;
	    RECT 105.1000 8.6000 105.4000 8.9000 ;
	    RECT 105.1000 8.3000 106.5000 8.6000 ;
	    RECT 106.1000 8.2000 106.5000 8.3000 ;
	    RECT 107.0000 7.8000 107.4000 8.6000 ;
	    RECT 107.8000 8.5000 108.2000 8.9000 ;
	    RECT 102.1000 7.7000 102.5000 7.8000 ;
	    RECT 94.2000 7.3000 95.3000 7.6000 ;
	    RECT 96.6000 7.3000 97.7000 7.6000 ;
	    RECT 94.2000 6.1000 94.6000 6.6000 ;
	    RECT 93.4000 5.8000 94.6000 6.1000 ;
	    RECT 95.0000 5.8000 95.3000 7.3000 ;
	    RECT 96.6000 5.8000 97.0000 6.6000 ;
	    RECT 97.4000 5.8000 97.7000 7.3000 ;
	    RECT 100.6000 7.4000 102.5000 7.7000 ;
	    RECT 76.6000 5.5000 79.4000 5.6000 ;
	    RECT 76.5000 5.4000 79.4000 5.5000 ;
	    RECT 80.4000 5.4000 81.0000 5.8000 ;
	    RECT 82.8000 5.4000 83.4000 5.8000 ;
	    RECT 72.6000 4.9000 73.8000 5.2000 ;
	    RECT 74.5000 5.3000 79.4000 5.4000 ;
	    RECT 74.5000 5.1000 76.9000 5.3000 ;
	    RECT 72.6000 4.4000 72.9000 4.9000 ;
	    RECT 72.2000 4.0000 72.9000 4.4000 ;
	    RECT 73.7000 4.5000 74.1000 4.6000 ;
	    RECT 74.5000 4.5000 74.8000 5.1000 ;
	    RECT 73.7000 4.2000 74.8000 4.5000 ;
	    RECT 75.1000 4.5000 77.8000 4.8000 ;
	    RECT 75.1000 4.4000 75.5000 4.5000 ;
	    RECT 77.4000 4.4000 77.8000 4.5000 ;
	    RECT 74.3000 3.7000 74.7000 3.8000 ;
	    RECT 75.7000 3.7000 76.1000 3.8000 ;
	    RECT 72.6000 3.1000 73.0000 3.5000 ;
	    RECT 74.3000 3.4000 76.1000 3.7000 ;
	    RECT 74.7000 3.1000 75.0000 3.4000 ;
	    RECT 77.4000 3.1000 77.8000 3.5000 ;
	    RECT 72.3000 1.1000 72.9000 3.1000 ;
	    RECT 74.6000 1.1000 75.0000 3.1000 ;
	    RECT 76.8000 2.8000 77.8000 3.1000 ;
	    RECT 76.8000 1.1000 77.2000 2.8000 ;
	    RECT 79.0000 1.1000 79.4000 5.3000 ;
	    RECT 80.7000 5.1000 81.0000 5.4000 ;
	    RECT 83.1000 5.1000 83.4000 5.4000 ;
	    RECT 84.6000 5.5000 87.4000 5.6000 ;
	    RECT 84.6000 5.4000 87.5000 5.5000 ;
	    RECT 84.6000 5.3000 89.5000 5.4000 ;
	    RECT 80.7000 4.8000 81.8000 5.1000 ;
	    RECT 83.1000 4.8000 84.2000 5.1000 ;
	    RECT 81.4000 1.1000 81.8000 4.8000 ;
	    RECT 83.8000 1.1000 84.2000 4.8000 ;
	    RECT 84.6000 1.1000 85.0000 5.3000 ;
	    RECT 87.1000 5.1000 89.5000 5.3000 ;
	    RECT 86.2000 4.5000 88.9000 4.8000 ;
	    RECT 86.2000 4.4000 86.6000 4.5000 ;
	    RECT 88.5000 4.4000 88.9000 4.5000 ;
	    RECT 89.2000 4.5000 89.5000 5.1000 ;
	    RECT 90.2000 5.2000 90.5000 5.8000 ;
	    RECT 91.7000 5.7000 92.1000 5.8000 ;
	    RECT 93.4000 5.7000 93.8000 5.8000 ;
	    RECT 91.7000 5.4000 93.8000 5.7000 ;
	    RECT 90.2000 4.9000 91.4000 5.2000 ;
	    RECT 89.9000 4.5000 90.3000 4.6000 ;
	    RECT 89.2000 4.2000 90.3000 4.5000 ;
	    RECT 91.1000 4.4000 91.4000 4.9000 ;
	    RECT 91.1000 4.0000 91.8000 4.4000 ;
	    RECT 87.9000 3.7000 88.3000 3.8000 ;
	    RECT 89.3000 3.7000 89.7000 3.8000 ;
	    RECT 86.2000 3.1000 86.6000 3.5000 ;
	    RECT 87.9000 3.4000 89.7000 3.7000 ;
	    RECT 89.0000 3.1000 89.3000 3.4000 ;
	    RECT 91.0000 3.1000 91.4000 3.5000 ;
	    RECT 86.2000 2.8000 87.2000 3.1000 ;
	    RECT 86.8000 1.1000 87.2000 2.8000 ;
	    RECT 89.0000 1.1000 89.4000 3.1000 ;
	    RECT 91.1000 1.1000 91.7000 3.1000 ;
	    RECT 93.4000 1.1000 93.8000 5.4000 ;
	    RECT 95.0000 5.4000 95.6000 5.8000 ;
	    RECT 97.4000 5.4000 98.0000 5.8000 ;
	    RECT 100.6000 5.7000 101.0000 7.4000 ;
	    RECT 104.1000 7.1000 104.5000 7.2000 ;
	    RECT 107.0000 7.1000 107.3000 7.8000 ;
	    RECT 109.4000 7.5000 109.8000 9.9000 ;
	    RECT 110.2000 7.6000 110.6000 9.9000 ;
	    RECT 112.6000 7.6000 113.0000 9.9000 ;
	    RECT 115.0000 7.6000 115.4000 9.9000 ;
	    RECT 110.2000 7.3000 111.3000 7.6000 ;
	    RECT 112.6000 7.3000 113.7000 7.6000 ;
	    RECT 115.0000 7.3000 116.1000 7.6000 ;
	    RECT 108.6000 7.1000 109.4000 7.2000 ;
	    RECT 103.9000 6.8000 109.4000 7.1000 ;
	    RECT 103.0000 6.4000 103.4000 6.5000 ;
	    RECT 101.5000 6.1000 103.4000 6.4000 ;
	    RECT 103.9000 6.1000 104.2000 6.8000 ;
	    RECT 107.5000 6.7000 107.9000 6.8000 ;
	    RECT 107.0000 6.2000 107.4000 6.3000 ;
	    RECT 108.3000 6.2000 108.7000 6.3000 ;
	    RECT 104.6000 6.1000 105.0000 6.2000 ;
	    RECT 101.5000 6.0000 101.9000 6.1000 ;
	    RECT 103.8000 5.8000 105.0000 6.1000 ;
	    RECT 106.2000 5.9000 108.7000 6.2000 ;
	    RECT 106.2000 5.8000 106.6000 5.9000 ;
	    RECT 110.2000 5.8000 110.6000 6.6000 ;
	    RECT 111.0000 5.8000 111.3000 7.3000 ;
	    RECT 112.6000 5.8000 113.0000 6.6000 ;
	    RECT 113.4000 5.8000 113.7000 7.3000 ;
	    RECT 115.0000 5.8000 115.4000 6.6000 ;
	    RECT 115.8000 5.8000 116.1000 7.3000 ;
	    RECT 116.6000 6.2000 117.0000 9.9000 ;
	    RECT 117.4000 7.6000 117.8000 9.9000 ;
	    RECT 117.4000 7.3000 118.5000 7.6000 ;
	    RECT 102.3000 5.7000 102.7000 5.8000 ;
	    RECT 100.6000 5.4000 102.7000 5.7000 ;
	    RECT 95.0000 5.1000 95.3000 5.4000 ;
	    RECT 97.4000 5.1000 97.7000 5.4000 ;
	    RECT 94.2000 4.8000 95.3000 5.1000 ;
	    RECT 96.6000 4.8000 97.7000 5.1000 ;
	    RECT 94.2000 1.1000 94.6000 4.8000 ;
	    RECT 96.6000 1.1000 97.0000 4.8000 ;
	    RECT 100.6000 1.1000 101.0000 5.4000 ;
	    RECT 103.9000 5.2000 104.2000 5.8000 ;
	    RECT 107.0000 5.5000 109.8000 5.6000 ;
	    RECT 106.9000 5.4000 109.8000 5.5000 ;
	    RECT 103.0000 4.9000 104.2000 5.2000 ;
	    RECT 104.9000 5.3000 109.8000 5.4000 ;
	    RECT 104.9000 5.1000 107.3000 5.3000 ;
	    RECT 103.0000 4.4000 103.3000 4.9000 ;
	    RECT 102.6000 4.0000 103.3000 4.4000 ;
	    RECT 104.1000 4.5000 104.5000 4.6000 ;
	    RECT 104.9000 4.5000 105.2000 5.1000 ;
	    RECT 104.1000 4.2000 105.2000 4.5000 ;
	    RECT 105.5000 4.5000 108.2000 4.8000 ;
	    RECT 105.5000 4.4000 105.9000 4.5000 ;
	    RECT 107.8000 4.4000 108.2000 4.5000 ;
	    RECT 104.7000 3.7000 105.1000 3.8000 ;
	    RECT 106.1000 3.7000 106.5000 3.8000 ;
	    RECT 103.0000 3.1000 103.4000 3.5000 ;
	    RECT 104.7000 3.4000 106.5000 3.7000 ;
	    RECT 105.1000 3.1000 105.4000 3.4000 ;
	    RECT 107.8000 3.1000 108.2000 3.5000 ;
	    RECT 102.7000 1.1000 103.3000 3.1000 ;
	    RECT 105.0000 1.1000 105.4000 3.1000 ;
	    RECT 107.2000 2.8000 108.2000 3.1000 ;
	    RECT 107.2000 1.1000 107.6000 2.8000 ;
	    RECT 109.4000 1.1000 109.8000 5.3000 ;
	    RECT 111.0000 5.4000 111.6000 5.8000 ;
	    RECT 113.4000 5.4000 114.0000 5.8000 ;
	    RECT 115.8000 5.4000 116.4000 5.8000 ;
	    RECT 111.0000 5.1000 111.3000 5.4000 ;
	    RECT 113.4000 5.1000 113.7000 5.4000 ;
	    RECT 115.8000 5.1000 116.1000 5.4000 ;
	    RECT 116.7000 5.1000 117.0000 6.2000 ;
	    RECT 117.4000 5.8000 117.8000 6.6000 ;
	    RECT 118.2000 5.8000 118.5000 7.3000 ;
	    RECT 119.0000 6.2000 119.4000 9.9000 ;
	    RECT 119.8000 7.6000 120.2000 9.9000 ;
	    RECT 122.2000 7.6000 122.6000 9.9000 ;
	    RECT 119.8000 7.3000 120.9000 7.6000 ;
	    RECT 122.2000 7.3000 123.3000 7.6000 ;
	    RECT 118.2000 5.4000 118.8000 5.8000 ;
	    RECT 118.2000 5.1000 118.5000 5.4000 ;
	    RECT 119.1000 5.1000 119.4000 6.2000 ;
	    RECT 119.8000 5.8000 120.2000 6.6000 ;
	    RECT 120.6000 5.8000 120.9000 7.3000 ;
	    RECT 122.2000 5.8000 122.6000 6.6000 ;
	    RECT 123.0000 5.8000 123.3000 7.3000 ;
	    RECT 123.8000 6.2000 124.2000 9.9000 ;
	    RECT 124.6000 7.6000 125.0000 9.9000 ;
	    RECT 127.0000 7.9000 127.4000 9.9000 ;
	    RECT 129.2000 9.2000 130.0000 9.9000 ;
	    RECT 129.2000 8.8000 130.6000 9.2000 ;
	    RECT 129.2000 8.1000 130.0000 8.8000 ;
	    RECT 127.0000 7.6000 128.3000 7.9000 ;
	    RECT 124.6000 7.3000 125.7000 7.6000 ;
	    RECT 127.9000 7.5000 128.3000 7.6000 ;
	    RECT 128.6000 7.4000 129.4000 7.8000 ;
	    RECT 120.6000 5.4000 121.2000 5.8000 ;
	    RECT 123.0000 5.4000 123.6000 5.8000 ;
	    RECT 120.6000 5.1000 120.9000 5.4000 ;
	    RECT 123.0000 5.1000 123.3000 5.4000 ;
	    RECT 123.9000 5.1000 124.2000 6.2000 ;
	    RECT 124.6000 5.8000 125.0000 6.6000 ;
	    RECT 125.4000 5.8000 125.7000 7.3000 ;
	    RECT 127.0000 7.1000 127.8000 7.2000 ;
	    RECT 129.7000 7.1000 130.0000 8.1000 ;
	    RECT 131.8000 7.9000 132.2000 9.9000 ;
	    RECT 130.3000 7.4000 130.7000 7.8000 ;
	    RECT 131.0000 7.6000 132.2000 7.9000 ;
	    RECT 132.6000 7.6000 133.0000 9.9000 ;
	    RECT 131.0000 7.5000 131.4000 7.6000 ;
	    RECT 127.0000 7.0000 128.1000 7.1000 ;
	    RECT 127.0000 6.8000 129.2000 7.0000 ;
	    RECT 127.8000 6.7000 129.2000 6.8000 ;
	    RECT 128.8000 6.6000 129.2000 6.7000 ;
	    RECT 129.5000 6.8000 130.0000 7.1000 ;
	    RECT 130.4000 7.2000 130.7000 7.4000 ;
	    RECT 132.6000 7.3000 133.7000 7.6000 ;
	    RECT 130.4000 6.8000 130.8000 7.2000 ;
	    RECT 131.4000 6.8000 132.2000 7.2000 ;
	    RECT 129.5000 6.2000 129.8000 6.8000 ;
	    RECT 128.1000 6.1000 128.5000 6.2000 ;
	    RECT 128.1000 5.8000 128.9000 6.1000 ;
	    RECT 129.4000 5.8000 129.8000 6.2000 ;
	    RECT 131.8000 6.1000 132.1000 6.8000 ;
	    RECT 132.6000 6.1000 133.0000 6.6000 ;
	    RECT 131.8000 5.8000 133.0000 6.1000 ;
	    RECT 133.4000 5.8000 133.7000 7.3000 ;
	    RECT 135.0000 6.2000 135.4000 9.9000 ;
	    RECT 136.6000 7.6000 137.0000 9.9000 ;
	    RECT 135.9000 7.3000 137.0000 7.6000 ;
	    RECT 137.4000 7.6000 137.8000 9.9000 ;
	    RECT 139.8000 7.6000 140.2000 9.9000 ;
	    RECT 142.2000 7.6000 142.6000 9.9000 ;
	    RECT 145.9000 9.2000 146.3000 9.9000 ;
	    RECT 145.4000 8.8000 146.3000 9.2000 ;
	    RECT 145.9000 8.2000 146.3000 8.8000 ;
	    RECT 145.4000 7.9000 146.3000 8.2000 ;
	    RECT 137.4000 7.3000 138.5000 7.6000 ;
	    RECT 139.8000 7.3000 140.9000 7.6000 ;
	    RECT 142.2000 7.3000 143.3000 7.6000 ;
	    RECT 125.4000 5.4000 126.0000 5.8000 ;
	    RECT 128.5000 5.7000 128.9000 5.8000 ;
	    RECT 125.4000 5.1000 125.7000 5.4000 ;
	    RECT 129.5000 5.1000 129.8000 5.8000 ;
	    RECT 133.4000 5.4000 134.0000 5.8000 ;
	    RECT 133.4000 5.1000 133.7000 5.4000 ;
	    RECT 110.2000 4.8000 111.3000 5.1000 ;
	    RECT 112.6000 4.8000 113.7000 5.1000 ;
	    RECT 115.0000 4.8000 116.1000 5.1000 ;
	    RECT 110.2000 1.1000 110.6000 4.8000 ;
	    RECT 112.6000 1.1000 113.0000 4.8000 ;
	    RECT 115.0000 1.1000 115.4000 4.8000 ;
	    RECT 116.6000 1.1000 117.0000 5.1000 ;
	    RECT 117.4000 4.8000 118.5000 5.1000 ;
	    RECT 117.4000 1.1000 117.8000 4.8000 ;
	    RECT 119.0000 1.1000 119.4000 5.1000 ;
	    RECT 119.8000 4.8000 120.9000 5.1000 ;
	    RECT 122.2000 4.8000 123.3000 5.1000 ;
	    RECT 119.8000 1.1000 120.2000 4.8000 ;
	    RECT 122.2000 1.1000 122.6000 4.8000 ;
	    RECT 123.8000 1.1000 124.2000 5.1000 ;
	    RECT 124.6000 4.8000 125.7000 5.1000 ;
	    RECT 127.0000 4.8000 128.3000 5.1000 ;
	    RECT 124.6000 1.1000 125.0000 4.8000 ;
	    RECT 127.0000 1.1000 127.4000 4.8000 ;
	    RECT 127.9000 4.7000 128.3000 4.8000 ;
	    RECT 129.2000 1.1000 130.0000 5.1000 ;
	    RECT 131.0000 4.8000 132.2000 5.1000 ;
	    RECT 131.0000 4.7000 131.4000 4.8000 ;
	    RECT 131.8000 1.1000 132.2000 4.8000 ;
	    RECT 132.6000 4.8000 133.7000 5.1000 ;
	    RECT 135.0000 5.1000 135.3000 6.2000 ;
	    RECT 135.9000 5.8000 136.2000 7.3000 ;
	    RECT 136.6000 6.1000 137.0000 6.6000 ;
	    RECT 137.4000 6.1000 137.8000 6.6000 ;
	    RECT 136.6000 5.8000 137.8000 6.1000 ;
	    RECT 138.2000 5.8000 138.5000 7.3000 ;
	    RECT 139.8000 5.8000 140.2000 6.6000 ;
	    RECT 140.6000 5.8000 140.9000 7.3000 ;
	    RECT 142.2000 5.8000 142.6000 6.6000 ;
	    RECT 143.0000 5.8000 143.3000 7.3000 ;
	    RECT 144.6000 6.8000 145.0000 7.6000 ;
	    RECT 135.6000 5.4000 136.2000 5.8000 ;
	    RECT 135.9000 5.1000 136.2000 5.4000 ;
	    RECT 138.2000 5.4000 138.8000 5.8000 ;
	    RECT 140.6000 5.4000 141.2000 5.8000 ;
	    RECT 143.0000 5.4000 143.6000 5.8000 ;
	    RECT 138.2000 5.1000 138.5000 5.4000 ;
	    RECT 140.6000 5.1000 140.9000 5.4000 ;
	    RECT 143.0000 5.1000 143.3000 5.4000 ;
	    RECT 132.6000 1.1000 133.0000 4.8000 ;
	    RECT 135.0000 1.1000 135.4000 5.1000 ;
	    RECT 135.9000 4.8000 137.0000 5.1000 ;
	    RECT 136.6000 1.1000 137.0000 4.8000 ;
	    RECT 137.4000 4.8000 138.5000 5.1000 ;
	    RECT 139.8000 4.8000 140.9000 5.1000 ;
	    RECT 142.2000 4.8000 143.3000 5.1000 ;
	    RECT 137.4000 1.1000 137.8000 4.8000 ;
	    RECT 139.8000 1.1000 140.2000 4.8000 ;
	    RECT 142.2000 1.1000 142.6000 4.8000 ;
	    RECT 145.4000 1.1000 145.8000 7.9000 ;
         LAYER metal2 ;
	    RECT 0.6000 116.8000 1.0000 117.2000 ;
	    RECT 0.6000 113.2000 0.9000 116.8000 ;
	    RECT 0.6000 112.8000 1.0000 113.2000 ;
	    RECT 3.0000 112.1000 3.4000 117.9000 ;
	    RECT 7.0000 115.8000 7.4000 116.2000 ;
	    RECT 7.0000 115.1000 7.3000 115.8000 ;
	    RECT 7.0000 114.7000 7.4000 115.1000 ;
	    RECT 7.0000 112.8000 7.4000 113.2000 ;
	    RECT 5.4000 103.1000 5.8000 108.9000 ;
	    RECT 6.2000 107.8000 6.6000 108.2000 ;
	    RECT 6.2000 107.2000 6.5000 107.8000 ;
	    RECT 6.2000 106.8000 6.6000 107.2000 ;
	    RECT 7.0000 106.2000 7.3000 112.8000 ;
	    RECT 7.8000 112.1000 8.2000 117.9000 ;
	    RECT 19.8000 116.8000 20.2000 117.2000 ;
	    RECT 21.4000 117.1000 21.8000 117.2000 ;
	    RECT 22.2000 117.1000 22.6000 117.2000 ;
	    RECT 21.4000 116.8000 22.6000 117.1000 ;
	    RECT 13.4000 115.9000 13.8000 116.3000 ;
	    RECT 9.4000 113.1000 9.8000 115.9000 ;
	    RECT 13.4000 114.2000 13.7000 115.9000 ;
	    RECT 14.2000 115.8000 14.6000 116.2000 ;
	    RECT 16.7000 115.9000 17.1000 116.3000 ;
	    RECT 14.2000 115.2000 14.5000 115.8000 ;
	    RECT 14.2000 114.8000 14.6000 115.2000 ;
	    RECT 15.4000 114.2000 15.8000 114.3000 ;
	    RECT 12.6000 113.8000 13.0000 114.2000 ;
	    RECT 13.4000 113.9000 15.8000 114.2000 ;
	    RECT 12.6000 113.2000 12.9000 113.8000 ;
	    RECT 13.4000 113.5000 13.7000 113.9000 ;
	    RECT 14.1000 113.5000 14.5000 113.6000 ;
	    RECT 15.8000 113.5000 16.2000 113.6000 ;
	    RECT 16.8000 113.5000 17.1000 115.9000 ;
	    RECT 19.8000 115.2000 20.1000 116.8000 ;
	    RECT 17.4000 114.8000 17.8000 115.2000 ;
	    RECT 19.8000 114.8000 20.2000 115.2000 ;
	    RECT 17.4000 114.2000 17.7000 114.8000 ;
	    RECT 17.4000 113.8000 17.8000 114.2000 ;
	    RECT 12.6000 112.8000 13.0000 113.2000 ;
	    RECT 13.4000 113.1000 13.8000 113.5000 ;
	    RECT 14.1000 113.2000 16.2000 113.5000 ;
	    RECT 16.7000 113.1000 17.1000 113.5000 ;
	    RECT 17.4000 113.1000 17.8000 113.2000 ;
	    RECT 18.2000 113.1000 18.6000 113.2000 ;
	    RECT 17.4000 112.8000 18.6000 113.1000 ;
	    RECT 19.0000 112.8000 19.4000 113.2000 ;
	    RECT 19.0000 112.2000 19.3000 112.8000 ;
	    RECT 19.0000 111.8000 19.4000 112.2000 ;
	    RECT 24.6000 112.1000 25.0000 117.9000 ;
	    RECT 25.4000 114.8000 25.8000 115.2000 ;
	    RECT 7.0000 105.8000 7.4000 106.2000 ;
	    RECT 8.6000 106.1000 9.0000 106.2000 ;
	    RECT 9.4000 106.1000 9.8000 106.3000 ;
	    RECT 8.6000 105.9000 9.8000 106.1000 ;
	    RECT 8.6000 105.8000 9.7000 105.9000 ;
	    RECT 7.0000 97.2000 7.3000 105.8000 ;
	    RECT 10.2000 103.1000 10.6000 108.9000 ;
	    RECT 11.8000 105.1000 12.2000 107.9000 ;
	    RECT 12.6000 107.8000 13.0000 108.2000 ;
	    RECT 12.6000 107.2000 12.9000 107.8000 ;
	    RECT 12.6000 106.8000 13.0000 107.2000 ;
	    RECT 14.2000 106.8000 14.6000 107.2000 ;
	    RECT 19.8000 107.1000 20.2000 107.2000 ;
	    RECT 20.6000 107.1000 21.0000 107.2000 ;
	    RECT 19.8000 106.8000 21.0000 107.1000 ;
	    RECT 14.2000 106.2000 14.5000 106.8000 ;
	    RECT 14.2000 105.8000 14.6000 106.2000 ;
	    RECT 15.8000 105.8000 16.2000 106.2000 ;
	    RECT 2.2000 96.8000 2.6000 97.2000 ;
	    RECT 7.0000 96.8000 7.4000 97.2000 ;
	    RECT 2.2000 95.2000 2.5000 96.8000 ;
	    RECT 2.2000 94.8000 2.6000 95.2000 ;
	    RECT 6.2000 93.8000 6.6000 94.2000 ;
	    RECT 4.6000 88.8000 5.0000 89.2000 ;
	    RECT 4.6000 88.2000 4.9000 88.8000 ;
	    RECT 4.6000 87.8000 5.0000 88.2000 ;
	    RECT 5.4000 83.1000 5.8000 88.9000 ;
	    RECT 6.2000 87.2000 6.5000 93.8000 ;
	    RECT 7.8000 92.1000 8.2000 97.9000 ;
	    RECT 11.8000 94.7000 12.2000 95.1000 ;
	    RECT 9.4000 93.8000 9.8000 94.2000 ;
	    RECT 9.4000 88.2000 9.7000 93.8000 ;
	    RECT 11.8000 92.2000 12.1000 94.7000 ;
	    RECT 11.8000 91.8000 12.2000 92.2000 ;
	    RECT 12.6000 92.1000 13.0000 97.9000 ;
	    RECT 14.2000 97.1000 14.6000 97.2000 ;
	    RECT 15.0000 97.1000 15.4000 97.2000 ;
	    RECT 14.2000 96.8000 15.4000 97.1000 ;
	    RECT 13.4000 94.8000 13.8000 95.2000 ;
	    RECT 13.4000 94.2000 13.7000 94.8000 ;
	    RECT 13.4000 93.8000 13.8000 94.2000 ;
	    RECT 14.2000 93.1000 14.6000 95.9000 ;
	    RECT 14.2000 91.8000 14.6000 92.2000 ;
	    RECT 14.2000 89.2000 14.5000 91.8000 ;
	    RECT 15.8000 90.2000 16.1000 105.8000 ;
	    RECT 21.4000 103.1000 21.8000 108.9000 ;
	    RECT 25.4000 108.2000 25.7000 114.8000 ;
	    RECT 28.6000 114.7000 29.0000 115.1000 ;
	    RECT 28.6000 111.2000 28.9000 114.7000 ;
	    RECT 29.4000 112.1000 29.8000 117.9000 ;
	    RECT 31.8000 116.8000 32.2000 117.2000 ;
	    RECT 66.2000 116.8000 66.6000 117.2000 ;
	    RECT 31.0000 113.1000 31.4000 115.9000 ;
	    RECT 31.8000 114.2000 32.1000 116.8000 ;
	    RECT 32.6000 115.9000 33.0000 116.3000 ;
	    RECT 35.7000 115.9000 36.1000 116.3000 ;
	    RECT 32.6000 114.2000 32.9000 115.9000 ;
	    RECT 35.1000 114.9000 35.5000 115.3000 ;
	    RECT 35.1000 114.2000 35.4000 114.9000 ;
	    RECT 31.8000 113.8000 32.2000 114.2000 ;
	    RECT 32.6000 113.9000 35.4000 114.2000 ;
	    RECT 32.6000 113.5000 32.9000 113.9000 ;
	    RECT 33.3000 113.5000 33.7000 113.6000 ;
	    RECT 35.0000 113.5000 35.4000 113.6000 ;
	    RECT 35.8000 113.5000 36.1000 115.9000 ;
	    RECT 39.8000 116.1000 40.2000 116.2000 ;
	    RECT 40.6000 116.1000 41.0000 116.2000 ;
	    RECT 39.8000 115.8000 41.0000 116.1000 ;
	    RECT 42.2000 115.8000 42.6000 116.2000 ;
	    RECT 59.7000 115.9000 60.1000 116.3000 ;
	    RECT 63.0000 115.9000 63.4000 116.3000 ;
	    RECT 66.2000 116.2000 66.5000 116.8000 ;
	    RECT 38.2000 114.8000 38.6000 115.2000 ;
	    RECT 39.0000 115.1000 39.4000 115.2000 ;
	    RECT 39.8000 115.1000 40.2000 115.2000 ;
	    RECT 39.0000 114.8000 40.2000 115.1000 ;
	    RECT 40.6000 114.8000 41.0000 115.2000 ;
	    RECT 41.4000 114.8000 41.8000 115.2000 ;
	    RECT 38.2000 114.2000 38.5000 114.8000 ;
	    RECT 32.6000 113.1000 33.0000 113.5000 ;
	    RECT 33.3000 113.2000 36.1000 113.5000 ;
	    RECT 35.7000 113.1000 36.1000 113.2000 ;
	    RECT 36.6000 113.8000 37.0000 114.2000 ;
	    RECT 37.4000 113.8000 37.8000 114.2000 ;
	    RECT 38.2000 113.8000 38.6000 114.2000 ;
	    RECT 36.6000 113.2000 36.9000 113.8000 ;
	    RECT 36.6000 112.8000 37.0000 113.2000 ;
	    RECT 33.4000 111.8000 33.8000 112.2000 ;
	    RECT 33.4000 111.2000 33.7000 111.8000 ;
	    RECT 37.4000 111.2000 37.7000 113.8000 ;
	    RECT 28.6000 110.8000 29.0000 111.2000 ;
	    RECT 33.4000 110.8000 33.8000 111.2000 ;
	    RECT 37.4000 110.8000 37.8000 111.2000 ;
	    RECT 38.2000 109.2000 38.5000 113.8000 ;
	    RECT 40.6000 112.2000 40.9000 114.8000 ;
	    RECT 41.4000 114.2000 41.7000 114.8000 ;
	    RECT 41.4000 113.8000 41.8000 114.2000 ;
	    RECT 40.6000 111.8000 41.0000 112.2000 ;
	    RECT 42.2000 109.2000 42.5000 115.8000 ;
	    RECT 43.8000 114.8000 44.2000 115.2000 ;
	    RECT 46.2000 114.8000 46.6000 115.2000 ;
	    RECT 52.6000 115.1000 53.0000 115.2000 ;
	    RECT 53.4000 115.1000 53.8000 115.2000 ;
	    RECT 52.6000 114.8000 53.8000 115.1000 ;
	    RECT 43.8000 114.2000 44.1000 114.8000 ;
	    RECT 43.8000 113.8000 44.2000 114.2000 ;
	    RECT 45.4000 113.8000 45.8000 114.2000 ;
	    RECT 45.4000 113.2000 45.7000 113.8000 ;
	    RECT 43.0000 112.8000 43.4000 113.2000 ;
	    RECT 43.8000 113.1000 44.2000 113.2000 ;
	    RECT 44.6000 113.1000 45.0000 113.2000 ;
	    RECT 43.8000 112.8000 45.0000 113.1000 ;
	    RECT 45.4000 112.8000 45.8000 113.2000 ;
	    RECT 43.0000 111.2000 43.3000 112.8000 ;
	    RECT 43.0000 110.8000 43.4000 111.2000 ;
	    RECT 25.4000 107.8000 25.8000 108.2000 ;
	    RECT 23.0000 105.8000 23.4000 106.2000 ;
	    RECT 25.4000 105.9000 25.8000 106.3000 ;
	    RECT 17.4000 92.1000 17.8000 97.9000 ;
	    RECT 19.0000 96.8000 19.4000 97.2000 ;
	    RECT 18.2000 93.8000 18.6000 94.2000 ;
	    RECT 18.2000 93.2000 18.5000 93.8000 ;
	    RECT 18.2000 92.8000 18.6000 93.2000 ;
	    RECT 15.8000 89.8000 16.2000 90.2000 ;
	    RECT 9.4000 87.8000 9.8000 88.2000 ;
	    RECT 6.2000 86.8000 6.6000 87.2000 ;
	    RECT 6.2000 75.2000 6.5000 86.8000 ;
	    RECT 9.4000 85.9000 9.8000 86.3000 ;
	    RECT 9.4000 84.2000 9.7000 85.9000 ;
	    RECT 9.4000 83.8000 9.8000 84.2000 ;
	    RECT 10.2000 83.1000 10.6000 88.9000 ;
	    RECT 14.2000 88.8000 14.6000 89.2000 ;
	    RECT 11.8000 85.1000 12.2000 87.9000 ;
	    RECT 12.6000 87.8000 13.0000 88.2000 ;
	    RECT 12.6000 87.2000 12.9000 87.8000 ;
	    RECT 13.4000 87.5000 13.8000 87.9000 ;
	    RECT 14.1000 87.5000 16.2000 87.8000 ;
	    RECT 16.7000 87.5000 17.1000 87.9000 ;
	    RECT 12.6000 86.8000 13.0000 87.2000 ;
	    RECT 13.4000 87.1000 13.7000 87.5000 ;
	    RECT 14.1000 87.4000 14.5000 87.5000 ;
	    RECT 15.8000 87.4000 16.2000 87.5000 ;
	    RECT 13.4000 86.8000 15.8000 87.1000 ;
	    RECT 13.4000 85.1000 13.7000 86.8000 ;
	    RECT 15.4000 86.7000 15.8000 86.8000 ;
	    RECT 16.8000 85.1000 17.1000 87.5000 ;
	    RECT 13.4000 84.7000 13.8000 85.1000 ;
	    RECT 16.7000 84.7000 17.1000 85.1000 ;
	    RECT 17.4000 86.8000 17.8000 87.2000 ;
	    RECT 18.2000 86.8000 18.6000 87.2000 ;
	    RECT 17.4000 85.1000 17.7000 86.8000 ;
	    RECT 18.2000 86.2000 18.5000 86.8000 ;
	    RECT 19.0000 86.2000 19.3000 96.8000 ;
	    RECT 21.4000 95.8000 21.8000 96.2000 ;
	    RECT 21.4000 95.1000 21.7000 95.8000 ;
	    RECT 21.4000 94.7000 21.8000 95.1000 ;
	    RECT 22.2000 92.1000 22.6000 97.9000 ;
	    RECT 23.0000 94.2000 23.3000 105.8000 ;
	    RECT 25.4000 105.2000 25.7000 105.9000 ;
	    RECT 25.4000 104.8000 25.8000 105.2000 ;
	    RECT 26.2000 103.1000 26.6000 108.9000 ;
	    RECT 38.2000 108.8000 38.6000 109.2000 ;
	    RECT 42.2000 108.8000 42.6000 109.2000 ;
	    RECT 27.8000 105.1000 28.2000 107.9000 ;
	    RECT 28.6000 107.8000 29.0000 108.2000 ;
	    RECT 39.0000 108.1000 39.4000 108.2000 ;
	    RECT 39.8000 108.1000 40.2000 108.2000 ;
	    RECT 28.6000 107.2000 28.9000 107.8000 ;
	    RECT 29.4000 107.5000 29.8000 107.9000 ;
	    RECT 30.1000 107.5000 32.2000 107.8000 ;
	    RECT 32.7000 107.5000 33.1000 107.9000 ;
	    RECT 39.0000 107.8000 40.2000 108.1000 ;
	    RECT 28.6000 106.8000 29.0000 107.2000 ;
	    RECT 29.4000 107.1000 29.7000 107.5000 ;
	    RECT 30.1000 107.4000 30.5000 107.5000 ;
	    RECT 31.8000 107.4000 32.2000 107.5000 ;
	    RECT 29.4000 106.8000 31.8000 107.1000 ;
	    RECT 28.6000 105.8000 29.0000 106.2000 ;
	    RECT 28.6000 105.2000 28.9000 105.8000 ;
	    RECT 28.6000 104.8000 29.0000 105.2000 ;
	    RECT 29.4000 105.1000 29.7000 106.8000 ;
	    RECT 31.4000 106.7000 31.8000 106.8000 ;
	    RECT 32.8000 105.1000 33.1000 107.5000 ;
	    RECT 29.4000 104.7000 29.8000 105.1000 ;
	    RECT 32.7000 104.7000 33.1000 105.1000 ;
	    RECT 33.4000 106.8000 33.8000 107.2000 ;
	    RECT 37.4000 107.1000 37.8000 107.2000 ;
	    RECT 38.2000 107.1000 38.6000 107.2000 ;
	    RECT 37.4000 106.8000 38.6000 107.1000 ;
	    RECT 33.4000 104.2000 33.7000 106.8000 ;
	    RECT 33.4000 103.8000 33.8000 104.2000 ;
	    RECT 39.8000 97.2000 40.1000 107.8000 ;
	    RECT 41.4000 106.8000 41.8000 107.2000 ;
	    RECT 41.4000 106.2000 41.7000 106.8000 ;
	    RECT 43.0000 106.2000 43.3000 110.8000 ;
	    RECT 46.2000 108.2000 46.5000 114.8000 ;
	    RECT 54.2000 113.8000 54.6000 114.2000 ;
	    RECT 51.8000 111.8000 52.2000 112.2000 ;
	    RECT 52.6000 111.8000 53.0000 112.2000 ;
	    RECT 46.2000 107.8000 46.6000 108.2000 ;
	    RECT 51.0000 107.8000 51.4000 108.2000 ;
	    RECT 51.0000 107.2000 51.3000 107.8000 ;
	    RECT 51.8000 107.2000 52.1000 111.8000 ;
	    RECT 52.6000 108.2000 52.9000 111.8000 ;
	    RECT 54.2000 111.2000 54.5000 113.8000 ;
	    RECT 59.7000 113.5000 60.0000 115.9000 ;
	    RECT 61.0000 114.2000 61.4000 114.3000 ;
	    RECT 63.1000 114.2000 63.4000 115.9000 ;
	    RECT 63.8000 115.8000 64.2000 116.2000 ;
	    RECT 64.6000 116.1000 65.0000 116.2000 ;
	    RECT 65.4000 116.1000 65.8000 116.2000 ;
	    RECT 64.6000 115.8000 65.8000 116.1000 ;
	    RECT 66.2000 115.8000 66.6000 116.2000 ;
	    RECT 63.8000 115.2000 64.1000 115.8000 ;
	    RECT 63.8000 114.8000 64.2000 115.2000 ;
	    RECT 61.0000 113.9000 63.4000 114.2000 ;
	    RECT 60.6000 113.5000 61.0000 113.6000 ;
	    RECT 62.3000 113.5000 62.7000 113.6000 ;
	    RECT 63.1000 113.5000 63.4000 113.9000 ;
	    RECT 64.6000 114.2000 64.9000 115.8000 ;
	    RECT 68.6000 114.8000 69.0000 115.2000 ;
	    RECT 64.6000 113.8000 65.0000 114.2000 ;
	    RECT 66.2000 113.8000 66.6000 114.2000 ;
	    RECT 67.8000 113.8000 68.2000 114.2000 ;
	    RECT 55.0000 112.8000 55.4000 113.2000 ;
	    RECT 55.8000 112.8000 56.2000 113.2000 ;
	    RECT 58.2000 112.8000 58.6000 113.2000 ;
	    RECT 59.7000 113.1000 60.1000 113.5000 ;
	    RECT 60.6000 113.2000 62.7000 113.5000 ;
	    RECT 63.0000 113.1000 63.4000 113.5000 ;
	    RECT 55.0000 112.2000 55.3000 112.8000 ;
	    RECT 55.0000 111.8000 55.4000 112.2000 ;
	    RECT 54.2000 110.8000 54.6000 111.2000 ;
	    RECT 55.8000 109.2000 56.1000 112.8000 ;
	    RECT 58.2000 112.2000 58.5000 112.8000 ;
	    RECT 58.2000 111.8000 58.6000 112.2000 ;
	    RECT 59.8000 111.8000 60.2000 112.2000 ;
	    RECT 64.6000 111.8000 65.0000 112.2000 ;
	    RECT 59.8000 109.2000 60.1000 111.8000 ;
	    RECT 63.0000 110.8000 63.4000 111.2000 ;
	    RECT 63.0000 109.2000 63.3000 110.8000 ;
	    RECT 55.8000 108.8000 56.2000 109.2000 ;
	    RECT 59.8000 108.8000 60.2000 109.2000 ;
	    RECT 63.0000 108.8000 63.4000 109.2000 ;
	    RECT 52.6000 107.8000 53.0000 108.2000 ;
	    RECT 47.0000 106.8000 47.4000 107.2000 ;
	    RECT 50.2000 106.8000 50.6000 107.2000 ;
	    RECT 51.0000 106.8000 51.4000 107.2000 ;
	    RECT 51.8000 106.8000 52.2000 107.2000 ;
	    RECT 55.0000 107.1000 55.4000 107.2000 ;
	    RECT 55.8000 107.1000 56.2000 107.2000 ;
	    RECT 55.0000 106.8000 56.2000 107.1000 ;
	    RECT 58.2000 107.1000 58.6000 107.2000 ;
	    RECT 59.0000 107.1000 59.4000 107.2000 ;
	    RECT 58.2000 106.8000 59.4000 107.1000 ;
	    RECT 61.4000 107.1000 61.8000 107.2000 ;
	    RECT 62.2000 107.1000 62.6000 107.2000 ;
	    RECT 61.4000 106.8000 62.6000 107.1000 ;
	    RECT 47.0000 106.2000 47.3000 106.8000 ;
	    RECT 50.2000 106.2000 50.5000 106.8000 ;
	    RECT 40.6000 105.8000 41.0000 106.2000 ;
	    RECT 41.4000 105.8000 41.8000 106.2000 ;
	    RECT 43.0000 105.8000 43.4000 106.2000 ;
	    RECT 43.8000 105.8000 44.2000 106.2000 ;
	    RECT 45.4000 105.8000 45.8000 106.2000 ;
	    RECT 47.0000 105.8000 47.4000 106.2000 ;
	    RECT 50.2000 105.8000 50.6000 106.2000 ;
	    RECT 58.2000 106.1000 58.6000 106.2000 ;
	    RECT 59.0000 106.1000 59.4000 106.2000 ;
	    RECT 58.2000 105.8000 59.4000 106.1000 ;
	    RECT 62.2000 105.8000 62.6000 106.2000 ;
	    RECT 24.6000 96.8000 25.0000 97.2000 ;
	    RECT 39.8000 96.8000 40.2000 97.2000 ;
	    RECT 23.0000 93.8000 23.4000 94.2000 ;
	    RECT 23.0000 89.2000 23.3000 93.8000 ;
	    RECT 23.8000 93.1000 24.2000 95.9000 ;
	    RECT 24.6000 94.2000 24.9000 96.8000 ;
	    RECT 25.4000 95.9000 25.8000 96.3000 ;
	    RECT 25.4000 94.2000 25.7000 95.9000 ;
	    RECT 26.2000 95.8000 26.6000 96.2000 ;
	    RECT 28.7000 95.9000 29.1000 96.3000 ;
	    RECT 26.2000 95.2000 26.5000 95.8000 ;
	    RECT 26.2000 94.8000 26.6000 95.2000 ;
	    RECT 27.4000 94.2000 27.8000 94.3000 ;
	    RECT 24.6000 93.8000 25.0000 94.2000 ;
	    RECT 25.4000 93.9000 27.8000 94.2000 ;
	    RECT 25.4000 93.5000 25.7000 93.9000 ;
	    RECT 26.1000 93.5000 26.5000 93.6000 ;
	    RECT 27.8000 93.5000 28.2000 93.6000 ;
	    RECT 28.8000 93.5000 29.1000 95.9000 ;
	    RECT 31.8000 96.1000 32.2000 96.2000 ;
	    RECT 32.6000 96.1000 33.0000 96.2000 ;
	    RECT 31.8000 95.8000 33.0000 96.1000 ;
	    RECT 36.6000 95.9000 37.0000 96.3000 ;
	    RECT 39.7000 95.9000 40.1000 96.3000 ;
	    RECT 29.4000 94.8000 29.8000 95.2000 ;
	    RECT 31.0000 95.1000 31.4000 95.2000 ;
	    RECT 31.8000 95.1000 32.2000 95.2000 ;
	    RECT 31.0000 94.8000 32.2000 95.1000 ;
	    RECT 32.6000 95.1000 33.0000 95.2000 ;
	    RECT 33.4000 95.1000 33.8000 95.2000 ;
	    RECT 32.6000 94.8000 33.8000 95.1000 ;
	    RECT 35.0000 95.1000 35.4000 95.2000 ;
	    RECT 35.8000 95.1000 36.2000 95.2000 ;
	    RECT 35.0000 94.8000 36.2000 95.1000 ;
	    RECT 29.4000 94.2000 29.7000 94.8000 ;
	    RECT 36.6000 94.2000 36.9000 95.9000 ;
	    RECT 39.1000 94.9000 39.5000 95.3000 ;
	    RECT 39.1000 94.2000 39.4000 94.9000 ;
	    RECT 29.4000 93.8000 29.8000 94.2000 ;
	    RECT 30.2000 93.8000 30.6000 94.2000 ;
	    RECT 31.8000 94.1000 32.2000 94.2000 ;
	    RECT 32.6000 94.1000 33.0000 94.2000 ;
	    RECT 31.8000 93.8000 33.0000 94.1000 ;
	    RECT 35.8000 93.8000 36.2000 94.2000 ;
	    RECT 36.6000 93.9000 39.4000 94.2000 ;
	    RECT 25.4000 93.1000 25.8000 93.5000 ;
	    RECT 26.1000 93.2000 28.2000 93.5000 ;
	    RECT 28.7000 93.1000 29.1000 93.5000 ;
	    RECT 30.2000 92.2000 30.5000 93.8000 ;
	    RECT 35.8000 93.2000 36.1000 93.8000 ;
	    RECT 36.6000 93.5000 36.9000 93.9000 ;
	    RECT 37.3000 93.5000 37.7000 93.6000 ;
	    RECT 39.0000 93.5000 39.4000 93.6000 ;
	    RECT 39.8000 93.5000 40.1000 95.9000 ;
	    RECT 40.6000 95.2000 40.9000 105.8000 ;
	    RECT 43.8000 105.2000 44.1000 105.8000 ;
	    RECT 45.4000 105.2000 45.7000 105.8000 ;
	    RECT 43.8000 104.8000 44.2000 105.2000 ;
	    RECT 45.4000 104.8000 45.8000 105.2000 ;
	    RECT 43.0000 96.8000 43.4000 97.2000 ;
	    RECT 40.6000 94.8000 41.0000 95.2000 ;
	    RECT 41.4000 94.8000 41.8000 95.2000 ;
	    RECT 33.4000 92.8000 33.8000 93.2000 ;
	    RECT 35.8000 92.8000 36.2000 93.2000 ;
	    RECT 36.6000 93.1000 37.0000 93.5000 ;
	    RECT 37.3000 93.2000 40.1000 93.5000 ;
	    RECT 39.7000 93.1000 40.1000 93.2000 ;
	    RECT 40.6000 93.8000 41.0000 94.2000 ;
	    RECT 40.6000 93.2000 40.9000 93.8000 ;
	    RECT 40.6000 92.8000 41.0000 93.2000 ;
	    RECT 27.0000 91.8000 27.4000 92.2000 ;
	    RECT 30.2000 91.8000 30.6000 92.2000 ;
	    RECT 24.6000 90.8000 25.0000 91.2000 ;
	    RECT 23.0000 88.8000 23.4000 89.2000 ;
	    RECT 23.0000 87.2000 23.3000 88.8000 ;
	    RECT 24.6000 88.2000 24.9000 90.8000 ;
	    RECT 27.0000 89.2000 27.3000 91.8000 ;
	    RECT 33.4000 91.2000 33.7000 92.8000 ;
	    RECT 41.4000 92.2000 41.7000 94.8000 ;
	    RECT 43.0000 94.2000 43.3000 96.8000 ;
	    RECT 43.8000 96.2000 44.1000 104.8000 ;
	    RECT 44.6000 103.8000 45.0000 104.2000 ;
	    RECT 44.6000 99.2000 44.9000 103.8000 ;
	    RECT 44.6000 98.8000 45.0000 99.2000 ;
	    RECT 43.8000 95.8000 44.2000 96.2000 ;
	    RECT 45.4000 95.2000 45.7000 104.8000 ;
	    RECT 44.6000 95.1000 45.0000 95.2000 ;
	    RECT 45.4000 95.1000 45.8000 95.2000 ;
	    RECT 44.6000 94.8000 45.8000 95.1000 ;
	    RECT 50.2000 94.2000 50.5000 105.8000 ;
	    RECT 55.8000 105.1000 56.2000 105.2000 ;
	    RECT 55.0000 104.8000 56.2000 105.1000 ;
	    RECT 56.6000 104.8000 57.0000 105.2000 ;
	    RECT 59.0000 105.1000 59.4000 105.2000 ;
	    RECT 59.8000 105.1000 60.2000 105.2000 ;
	    RECT 59.0000 104.8000 60.2000 105.1000 ;
	    RECT 55.0000 99.2000 55.3000 104.8000 ;
	    RECT 55.0000 98.8000 55.4000 99.2000 ;
	    RECT 56.6000 96.2000 56.9000 104.8000 ;
	    RECT 58.2000 97.1000 58.6000 97.2000 ;
	    RECT 59.0000 97.1000 59.4000 97.2000 ;
	    RECT 58.2000 96.8000 59.4000 97.1000 ;
	    RECT 56.6000 95.8000 57.0000 96.2000 ;
	    RECT 57.4000 95.8000 57.8000 96.2000 ;
	    RECT 51.0000 94.8000 51.4000 95.2000 ;
	    RECT 54.2000 95.1000 54.6000 95.2000 ;
	    RECT 55.0000 95.1000 55.4000 95.2000 ;
	    RECT 54.2000 94.8000 55.4000 95.1000 ;
	    RECT 43.0000 93.8000 43.4000 94.2000 ;
	    RECT 50.2000 94.1000 50.6000 94.2000 ;
	    RECT 49.4000 93.8000 50.6000 94.1000 ;
	    RECT 43.0000 93.2000 43.3000 93.8000 ;
	    RECT 43.0000 92.8000 43.4000 93.2000 ;
	    RECT 48.6000 92.8000 49.0000 93.2000 ;
	    RECT 37.4000 91.8000 37.8000 92.2000 ;
	    RECT 41.4000 91.8000 41.8000 92.2000 ;
	    RECT 33.4000 90.8000 33.8000 91.2000 ;
	    RECT 27.0000 88.8000 27.4000 89.2000 ;
	    RECT 28.6000 88.8000 29.0000 89.2000 ;
	    RECT 24.6000 87.8000 25.0000 88.2000 ;
	    RECT 27.8000 87.8000 28.2000 88.2000 ;
	    RECT 23.0000 86.8000 23.4000 87.2000 ;
	    RECT 24.6000 86.2000 24.9000 87.8000 ;
	    RECT 18.2000 85.8000 18.6000 86.2000 ;
	    RECT 19.0000 85.8000 19.4000 86.2000 ;
	    RECT 24.6000 85.8000 25.0000 86.2000 ;
	    RECT 17.4000 84.8000 18.5000 85.1000 ;
	    RECT 13.4000 82.8000 13.8000 83.2000 ;
	    RECT 12.6000 76.8000 13.0000 77.2000 ;
	    RECT 12.6000 76.2000 12.9000 76.8000 ;
	    RECT 12.6000 75.8000 13.0000 76.2000 ;
	    RECT 13.4000 75.2000 13.7000 82.8000 ;
	    RECT 18.2000 79.2000 18.5000 84.8000 ;
	    RECT 19.0000 83.2000 19.3000 85.8000 ;
	    RECT 27.8000 85.2000 28.1000 87.8000 ;
	    RECT 28.6000 87.2000 28.9000 88.8000 ;
	    RECT 29.4000 87.5000 29.8000 87.9000 ;
	    RECT 30.1000 87.5000 32.2000 87.8000 ;
	    RECT 32.7000 87.5000 33.1000 87.9000 ;
	    RECT 28.6000 86.8000 29.0000 87.2000 ;
	    RECT 29.4000 87.1000 29.7000 87.5000 ;
	    RECT 30.1000 87.4000 30.5000 87.5000 ;
	    RECT 31.8000 87.4000 32.2000 87.5000 ;
	    RECT 29.4000 86.8000 31.8000 87.1000 ;
	    RECT 20.6000 85.1000 21.0000 85.2000 ;
	    RECT 21.4000 85.1000 21.8000 85.2000 ;
	    RECT 20.6000 84.8000 21.8000 85.1000 ;
	    RECT 27.8000 84.8000 28.2000 85.2000 ;
	    RECT 29.4000 85.1000 29.7000 86.8000 ;
	    RECT 31.4000 86.7000 31.8000 86.8000 ;
	    RECT 32.8000 85.1000 33.1000 87.5000 ;
	    RECT 33.4000 86.8000 33.8000 87.2000 ;
	    RECT 33.4000 86.2000 33.7000 86.8000 ;
	    RECT 33.4000 85.8000 33.8000 86.2000 ;
	    RECT 34.2000 85.1000 34.6000 87.9000 ;
	    RECT 35.0000 87.8000 35.4000 88.2000 ;
	    RECT 35.0000 87.2000 35.3000 87.8000 ;
	    RECT 35.0000 86.8000 35.4000 87.2000 ;
	    RECT 19.0000 82.8000 19.4000 83.2000 ;
	    RECT 19.0000 81.8000 19.4000 82.2000 ;
	    RECT 18.2000 78.8000 18.6000 79.2000 ;
	    RECT 15.8000 76.8000 16.2000 77.2000 ;
	    RECT 15.8000 76.2000 16.1000 76.8000 ;
	    RECT 15.8000 75.8000 16.2000 76.2000 ;
	    RECT 16.6000 76.1000 17.0000 76.2000 ;
	    RECT 17.4000 76.1000 17.8000 76.2000 ;
	    RECT 16.6000 75.8000 17.8000 76.1000 ;
	    RECT 19.0000 75.2000 19.3000 81.8000 ;
	    RECT 27.8000 79.2000 28.1000 84.8000 ;
	    RECT 29.4000 84.7000 29.8000 85.1000 ;
	    RECT 32.7000 84.7000 33.1000 85.1000 ;
	    RECT 30.2000 84.1000 30.6000 84.2000 ;
	    RECT 31.0000 84.1000 31.4000 84.2000 ;
	    RECT 30.2000 83.8000 31.4000 84.1000 ;
	    RECT 34.2000 83.8000 34.6000 84.2000 ;
	    RECT 34.2000 79.2000 34.5000 83.8000 ;
	    RECT 35.8000 83.1000 36.2000 88.9000 ;
	    RECT 37.4000 86.2000 37.7000 91.8000 ;
	    RECT 43.0000 89.2000 43.3000 92.8000 ;
	    RECT 37.4000 85.8000 37.8000 86.2000 ;
	    RECT 40.6000 83.1000 41.0000 88.9000 ;
	    RECT 43.0000 88.8000 43.4000 89.2000 ;
	    RECT 46.2000 88.8000 46.6000 89.2000 ;
	    RECT 43.0000 86.2000 43.3000 88.8000 ;
	    RECT 43.0000 85.8000 43.4000 86.2000 ;
	    RECT 44.6000 86.1000 45.0000 86.2000 ;
	    RECT 45.4000 86.1000 45.8000 86.2000 ;
	    RECT 44.6000 85.8000 45.8000 86.1000 ;
	    RECT 46.2000 85.2000 46.5000 88.8000 ;
	    RECT 47.0000 87.1000 47.4000 87.2000 ;
	    RECT 47.8000 87.1000 48.2000 87.2000 ;
	    RECT 47.0000 86.8000 48.2000 87.1000 ;
	    RECT 48.6000 86.2000 48.9000 92.8000 ;
	    RECT 48.6000 85.8000 49.0000 86.2000 ;
	    RECT 49.4000 85.2000 49.7000 93.8000 ;
	    RECT 51.0000 93.1000 51.3000 94.8000 ;
	    RECT 52.6000 93.8000 53.0000 94.2000 ;
	    RECT 53.4000 93.8000 53.8000 94.2000 ;
	    RECT 52.6000 93.2000 52.9000 93.8000 ;
	    RECT 50.2000 92.8000 51.3000 93.1000 ;
	    RECT 51.8000 92.8000 52.2000 93.2000 ;
	    RECT 52.6000 92.8000 53.0000 93.2000 ;
	    RECT 50.2000 86.2000 50.5000 92.8000 ;
	    RECT 51.8000 89.2000 52.1000 92.8000 ;
	    RECT 53.4000 92.2000 53.7000 93.8000 ;
	    RECT 53.4000 91.8000 53.8000 92.2000 ;
	    RECT 51.8000 88.8000 52.2000 89.2000 ;
	    RECT 53.4000 88.8000 53.8000 89.2000 ;
	    RECT 51.0000 87.8000 51.4000 88.2000 ;
	    RECT 51.0000 87.2000 51.3000 87.8000 ;
	    RECT 51.0000 86.8000 51.4000 87.2000 ;
	    RECT 53.4000 86.2000 53.7000 88.8000 ;
	    RECT 54.2000 87.2000 54.5000 94.8000 ;
	    RECT 55.8000 93.8000 56.2000 94.2000 ;
	    RECT 55.8000 93.2000 56.1000 93.8000 ;
	    RECT 55.8000 92.8000 56.2000 93.2000 ;
	    RECT 56.6000 92.1000 56.9000 95.8000 ;
	    RECT 57.4000 95.2000 57.7000 95.8000 ;
	    RECT 62.2000 95.2000 62.5000 105.8000 ;
	    RECT 64.6000 105.2000 64.9000 111.8000 ;
	    RECT 65.4000 106.8000 65.8000 107.2000 ;
	    RECT 65.4000 106.2000 65.7000 106.8000 ;
	    RECT 65.4000 105.8000 65.8000 106.2000 ;
	    RECT 63.0000 105.1000 63.4000 105.2000 ;
	    RECT 63.8000 105.1000 64.2000 105.2000 ;
	    RECT 63.0000 104.8000 64.2000 105.1000 ;
	    RECT 64.6000 104.8000 65.0000 105.2000 ;
	    RECT 63.0000 96.2000 63.3000 104.8000 ;
	    RECT 65.4000 103.8000 65.8000 104.2000 ;
	    RECT 64.6000 96.8000 65.0000 97.2000 ;
	    RECT 64.6000 96.2000 64.9000 96.8000 ;
	    RECT 65.4000 96.2000 65.7000 103.8000 ;
	    RECT 63.0000 95.8000 63.4000 96.2000 ;
	    RECT 64.6000 95.8000 65.0000 96.2000 ;
	    RECT 65.4000 95.8000 65.8000 96.2000 ;
	    RECT 57.4000 94.8000 57.8000 95.2000 ;
	    RECT 59.8000 94.8000 60.2000 95.2000 ;
	    RECT 62.2000 94.8000 62.6000 95.2000 ;
	    RECT 63.0000 94.8000 63.4000 95.2000 ;
	    RECT 57.4000 93.8000 57.8000 94.2000 ;
	    RECT 57.4000 93.2000 57.7000 93.8000 ;
	    RECT 57.4000 92.8000 57.8000 93.2000 ;
	    RECT 55.8000 91.8000 56.9000 92.1000 ;
	    RECT 58.2000 91.8000 58.6000 92.2000 ;
	    RECT 55.8000 87.2000 56.1000 91.8000 ;
	    RECT 58.2000 89.2000 58.5000 91.8000 ;
	    RECT 56.6000 88.8000 57.0000 89.2000 ;
	    RECT 58.2000 88.8000 58.6000 89.2000 ;
	    RECT 56.6000 88.2000 56.9000 88.8000 ;
	    RECT 59.8000 88.2000 60.1000 94.8000 ;
	    RECT 62.2000 93.2000 62.5000 94.8000 ;
	    RECT 63.0000 94.2000 63.3000 94.8000 ;
	    RECT 63.0000 93.8000 63.4000 94.2000 ;
	    RECT 62.2000 92.8000 62.6000 93.2000 ;
	    RECT 61.4000 89.1000 61.8000 89.2000 ;
	    RECT 62.2000 89.1000 62.6000 89.2000 ;
	    RECT 61.4000 88.8000 62.6000 89.1000 ;
	    RECT 56.6000 87.8000 57.0000 88.2000 ;
	    RECT 59.8000 87.8000 60.2000 88.2000 ;
	    RECT 64.6000 88.1000 65.0000 88.2000 ;
	    RECT 65.4000 88.1000 65.8000 88.2000 ;
	    RECT 64.6000 87.8000 65.8000 88.1000 ;
	    RECT 54.2000 86.8000 54.6000 87.2000 ;
	    RECT 55.8000 86.8000 56.2000 87.2000 ;
	    RECT 56.6000 86.8000 57.0000 87.2000 ;
	    RECT 57.4000 86.8000 57.8000 87.2000 ;
	    RECT 50.2000 85.8000 50.6000 86.2000 ;
	    RECT 51.0000 85.8000 51.4000 86.2000 ;
	    RECT 53.4000 85.8000 53.8000 86.2000 ;
	    RECT 54.2000 85.8000 54.6000 86.2000 ;
	    RECT 45.4000 84.8000 45.8000 85.2000 ;
	    RECT 46.2000 84.8000 46.6000 85.2000 ;
	    RECT 47.8000 84.8000 48.2000 85.2000 ;
	    RECT 49.4000 84.8000 49.8000 85.2000 ;
	    RECT 43.8000 84.1000 44.2000 84.2000 ;
	    RECT 44.6000 84.1000 45.0000 84.2000 ;
	    RECT 43.8000 83.8000 45.0000 84.1000 ;
	    RECT 45.4000 83.2000 45.7000 84.8000 ;
	    RECT 47.8000 83.2000 48.1000 84.8000 ;
	    RECT 43.8000 82.8000 44.2000 83.2000 ;
	    RECT 45.4000 82.8000 45.8000 83.2000 ;
	    RECT 47.8000 82.8000 48.2000 83.2000 ;
	    RECT 43.8000 79.2000 44.1000 82.8000 ;
	    RECT 27.8000 78.8000 28.2000 79.2000 ;
	    RECT 34.2000 78.8000 34.6000 79.2000 ;
	    RECT 43.8000 78.8000 44.2000 79.2000 ;
	    RECT 51.0000 78.2000 51.3000 85.8000 ;
	    RECT 51.8000 84.8000 52.2000 85.2000 ;
	    RECT 51.8000 83.2000 52.1000 84.8000 ;
	    RECT 53.4000 83.8000 53.8000 84.2000 ;
	    RECT 51.8000 82.8000 52.2000 83.2000 ;
	    RECT 53.4000 79.2000 53.7000 83.8000 ;
	    RECT 53.4000 78.8000 53.8000 79.2000 ;
	    RECT 35.8000 77.8000 36.2000 78.2000 ;
	    RECT 51.0000 77.8000 51.4000 78.2000 ;
	    RECT 24.6000 76.8000 25.0000 77.2000 ;
	    RECT 20.6000 75.8000 21.0000 76.2000 ;
	    RECT 3.8000 74.8000 4.2000 75.2000 ;
	    RECT 6.2000 74.8000 6.6000 75.2000 ;
	    RECT 7.0000 74.8000 7.4000 75.2000 ;
	    RECT 13.4000 74.8000 13.8000 75.2000 ;
	    RECT 19.0000 74.8000 19.4000 75.2000 ;
	    RECT 3.8000 73.2000 4.1000 74.8000 ;
	    RECT 7.0000 74.2000 7.3000 74.8000 ;
	    RECT 6.2000 73.8000 6.6000 74.2000 ;
	    RECT 7.0000 73.8000 7.4000 74.2000 ;
	    RECT 9.4000 73.8000 9.8000 74.2000 ;
	    RECT 10.2000 74.0000 10.6000 74.4000 ;
	    RECT 11.8000 74.1000 12.2000 74.2000 ;
	    RECT 12.6000 74.1000 13.0000 74.2000 ;
	    RECT 6.2000 73.2000 6.5000 73.8000 ;
	    RECT 9.4000 73.2000 9.7000 73.8000 ;
	    RECT 3.8000 72.8000 4.2000 73.2000 ;
	    RECT 5.4000 73.1000 5.8000 73.2000 ;
	    RECT 6.2000 73.1000 6.6000 73.2000 ;
	    RECT 5.4000 72.8000 6.6000 73.1000 ;
	    RECT 9.4000 72.8000 9.8000 73.2000 ;
	    RECT 3.8000 67.1000 4.2000 67.2000 ;
	    RECT 4.6000 67.1000 5.0000 67.2000 ;
	    RECT 3.8000 66.8000 5.0000 67.1000 ;
	    RECT 5.4000 63.1000 5.8000 68.9000 ;
	    RECT 6.2000 59.2000 6.5000 72.8000 ;
	    RECT 10.2000 72.2000 10.5000 74.0000 ;
	    RECT 11.8000 73.8000 13.0000 74.1000 ;
	    RECT 15.8000 73.8000 16.2000 74.2000 ;
	    RECT 15.8000 73.2000 16.1000 73.8000 ;
	    RECT 20.6000 73.2000 20.9000 75.8000 ;
	    RECT 24.6000 74.2000 24.9000 76.8000 ;
	    RECT 25.4000 76.1000 25.8000 76.2000 ;
	    RECT 26.2000 76.1000 26.6000 76.2000 ;
	    RECT 25.4000 75.8000 26.6000 76.1000 ;
	    RECT 31.0000 75.8000 31.4000 76.2000 ;
	    RECT 23.0000 74.1000 23.4000 74.2000 ;
	    RECT 23.8000 74.1000 24.2000 74.2000 ;
	    RECT 23.0000 73.8000 24.2000 74.1000 ;
	    RECT 24.6000 73.8000 25.0000 74.2000 ;
	    RECT 25.4000 73.2000 25.7000 75.8000 ;
	    RECT 31.0000 75.2000 31.3000 75.8000 ;
	    RECT 29.4000 75.1000 29.8000 75.2000 ;
	    RECT 30.2000 75.1000 30.6000 75.2000 ;
	    RECT 29.4000 74.8000 30.6000 75.1000 ;
	    RECT 31.0000 74.8000 31.4000 75.2000 ;
	    RECT 27.8000 73.8000 28.2000 74.2000 ;
	    RECT 27.8000 73.2000 28.1000 73.8000 ;
	    RECT 15.8000 72.8000 16.2000 73.2000 ;
	    RECT 20.6000 72.8000 21.0000 73.2000 ;
	    RECT 23.0000 72.8000 23.4000 73.2000 ;
	    RECT 23.8000 73.1000 24.2000 73.2000 ;
	    RECT 24.6000 73.1000 25.0000 73.2000 ;
	    RECT 23.8000 72.8000 25.0000 73.1000 ;
	    RECT 25.4000 72.8000 25.8000 73.2000 ;
	    RECT 27.8000 72.8000 28.2000 73.2000 ;
	    RECT 28.6000 72.8000 29.0000 73.2000 ;
	    RECT 29.4000 73.1000 29.8000 73.2000 ;
	    RECT 30.2000 73.1000 30.6000 73.2000 ;
	    RECT 29.4000 72.8000 30.6000 73.1000 ;
	    RECT 31.0000 72.8000 31.4000 73.2000 ;
	    RECT 32.6000 72.8000 33.0000 73.2000 ;
	    RECT 7.0000 71.8000 7.4000 72.2000 ;
	    RECT 10.2000 71.8000 10.6000 72.2000 ;
	    RECT 12.6000 71.8000 13.0000 72.2000 ;
	    RECT 17.4000 71.8000 17.8000 72.2000 ;
	    RECT 7.0000 69.2000 7.3000 71.8000 ;
	    RECT 7.0000 68.8000 7.4000 69.2000 ;
	    RECT 9.4000 65.9000 9.8000 66.3000 ;
	    RECT 9.4000 65.2000 9.7000 65.9000 ;
	    RECT 9.4000 64.8000 9.8000 65.2000 ;
	    RECT 10.2000 63.1000 10.6000 68.9000 ;
	    RECT 12.6000 68.2000 12.9000 71.8000 ;
	    RECT 17.4000 70.2000 17.7000 71.8000 ;
	    RECT 17.4000 69.8000 17.8000 70.2000 ;
	    RECT 20.6000 69.8000 21.0000 70.2000 ;
	    RECT 11.0000 66.8000 11.4000 67.2000 ;
	    RECT 6.2000 58.8000 6.6000 59.2000 ;
	    RECT 8.6000 59.1000 9.0000 59.2000 ;
	    RECT 9.4000 59.1000 9.8000 59.2000 ;
	    RECT 8.6000 58.8000 9.8000 59.1000 ;
	    RECT 11.0000 57.2000 11.3000 66.8000 ;
	    RECT 11.8000 65.1000 12.2000 67.9000 ;
	    RECT 12.6000 67.8000 13.0000 68.2000 ;
	    RECT 12.6000 67.2000 12.9000 67.8000 ;
	    RECT 15.0000 67.5000 15.4000 67.9000 ;
	    RECT 15.7000 67.5000 17.8000 67.8000 ;
	    RECT 18.3000 67.5000 18.7000 67.9000 ;
	    RECT 12.6000 66.8000 13.0000 67.2000 ;
	    RECT 14.2000 66.8000 14.6000 67.2000 ;
	    RECT 15.0000 67.1000 15.3000 67.5000 ;
	    RECT 15.7000 67.4000 16.1000 67.5000 ;
	    RECT 17.4000 67.4000 17.8000 67.5000 ;
	    RECT 15.0000 66.8000 17.4000 67.1000 ;
	    RECT 14.2000 66.2000 14.5000 66.8000 ;
	    RECT 14.2000 65.8000 14.6000 66.2000 ;
	    RECT 15.0000 65.1000 15.3000 66.8000 ;
	    RECT 17.0000 66.7000 17.4000 66.8000 ;
	    RECT 15.8000 65.8000 16.2000 66.2000 ;
	    RECT 15.8000 65.2000 16.1000 65.8000 ;
	    RECT 15.0000 64.7000 15.4000 65.1000 ;
	    RECT 15.8000 64.8000 16.2000 65.2000 ;
	    RECT 18.4000 65.1000 18.7000 67.5000 ;
	    RECT 19.0000 67.8000 19.4000 68.2000 ;
	    RECT 19.0000 67.2000 19.3000 67.8000 ;
	    RECT 20.6000 67.2000 20.9000 69.8000 ;
	    RECT 21.4000 68.1000 21.8000 68.2000 ;
	    RECT 22.2000 68.1000 22.6000 68.2000 ;
	    RECT 21.4000 67.8000 22.6000 68.1000 ;
	    RECT 19.0000 66.8000 19.4000 67.2000 ;
	    RECT 20.6000 66.8000 21.0000 67.2000 ;
	    RECT 19.8000 66.1000 20.2000 66.2000 ;
	    RECT 20.6000 66.1000 21.0000 66.2000 ;
	    RECT 19.8000 65.8000 21.0000 66.1000 ;
	    RECT 18.3000 64.7000 18.7000 65.1000 ;
	    RECT 23.0000 65.2000 23.3000 72.8000 ;
	    RECT 25.4000 72.1000 25.8000 72.2000 ;
	    RECT 26.2000 72.1000 26.6000 72.2000 ;
	    RECT 25.4000 71.8000 26.6000 72.1000 ;
	    RECT 25.4000 68.8000 25.8000 69.2000 ;
	    RECT 27.0000 68.8000 27.4000 69.2000 ;
	    RECT 25.4000 67.2000 25.7000 68.8000 ;
	    RECT 25.4000 66.8000 25.8000 67.2000 ;
	    RECT 24.6000 66.1000 25.0000 66.2000 ;
	    RECT 25.4000 66.1000 25.8000 66.2000 ;
	    RECT 24.6000 65.8000 25.8000 66.1000 ;
	    RECT 23.0000 65.1000 23.4000 65.2000 ;
	    RECT 23.0000 64.8000 24.1000 65.1000 ;
	    RECT 19.0000 58.8000 19.4000 59.2000 ;
	    RECT 11.0000 56.8000 11.4000 57.2000 ;
	    RECT 2.2000 54.8000 2.6000 55.2000 ;
	    RECT 4.6000 55.1000 5.0000 55.2000 ;
	    RECT 5.4000 55.1000 5.8000 55.2000 ;
	    RECT 4.6000 54.8000 5.8000 55.1000 ;
	    RECT 8.6000 55.1000 9.0000 55.2000 ;
	    RECT 9.4000 55.1000 9.8000 55.2000 ;
	    RECT 8.6000 54.8000 9.8000 55.1000 ;
	    RECT 2.2000 53.2000 2.5000 54.8000 ;
	    RECT 0.6000 52.8000 1.0000 53.2000 ;
	    RECT 2.2000 52.8000 2.6000 53.2000 ;
	    RECT 4.6000 53.1000 5.0000 53.2000 ;
	    RECT 5.4000 53.1000 5.8000 53.2000 ;
	    RECT 4.6000 52.8000 5.8000 53.1000 ;
	    RECT 0.6000 49.2000 0.9000 52.8000 ;
	    RECT 6.2000 51.8000 6.6000 52.2000 ;
	    RECT 11.8000 52.1000 12.2000 57.9000 ;
	    RECT 15.8000 55.8000 16.2000 56.2000 ;
	    RECT 12.6000 54.8000 13.0000 55.2000 ;
	    RECT 15.8000 55.1000 16.1000 55.8000 ;
	    RECT 6.2000 49.2000 6.5000 51.8000 ;
	    RECT 0.6000 48.8000 1.0000 49.2000 ;
	    RECT 3.0000 43.1000 3.4000 48.9000 ;
	    RECT 6.2000 48.8000 6.6000 49.2000 ;
	    RECT 7.0000 46.8000 7.4000 47.2000 ;
	    RECT 7.0000 46.3000 7.3000 46.8000 ;
	    RECT 7.0000 45.9000 7.4000 46.3000 ;
	    RECT 7.0000 45.8000 7.3000 45.9000 ;
	    RECT 7.8000 43.1000 8.2000 48.9000 ;
	    RECT 10.2000 48.8000 10.6000 49.2000 ;
	    RECT 10.2000 48.2000 10.5000 48.8000 ;
	    RECT 8.6000 47.8000 9.0000 48.2000 ;
	    RECT 8.6000 47.2000 8.9000 47.8000 ;
	    RECT 8.6000 46.8000 9.0000 47.2000 ;
	    RECT 5.4000 32.1000 5.8000 37.9000 ;
	    RECT 8.6000 34.2000 8.9000 46.8000 ;
	    RECT 9.4000 45.1000 9.8000 47.9000 ;
	    RECT 10.2000 47.8000 10.6000 48.2000 ;
	    RECT 10.2000 46.8000 10.6000 47.2000 ;
	    RECT 11.8000 46.8000 12.2000 47.2000 ;
	    RECT 10.2000 46.2000 10.5000 46.8000 ;
	    RECT 11.8000 46.2000 12.1000 46.8000 ;
	    RECT 12.6000 46.2000 12.9000 54.8000 ;
	    RECT 15.8000 54.7000 16.2000 55.1000 ;
	    RECT 16.6000 52.1000 17.0000 57.9000 ;
	    RECT 17.4000 53.8000 17.8000 54.2000 ;
	    RECT 17.4000 48.2000 17.7000 53.8000 ;
	    RECT 18.2000 53.1000 18.6000 55.9000 ;
	    RECT 19.0000 54.2000 19.3000 58.8000 ;
	    RECT 19.9000 55.9000 20.3000 56.3000 ;
	    RECT 23.0000 55.9000 23.4000 56.3000 ;
	    RECT 19.0000 53.8000 19.4000 54.2000 ;
	    RECT 19.9000 53.5000 20.2000 55.9000 ;
	    RECT 20.5000 54.9000 20.9000 55.3000 ;
	    RECT 20.6000 54.2000 20.9000 54.9000 ;
	    RECT 21.4000 55.1000 21.8000 55.2000 ;
	    RECT 22.2000 55.1000 22.6000 55.2000 ;
	    RECT 21.4000 54.8000 22.6000 55.1000 ;
	    RECT 23.1000 54.2000 23.4000 55.9000 ;
	    RECT 20.6000 53.9000 23.4000 54.2000 ;
	    RECT 20.6000 53.5000 21.0000 53.6000 ;
	    RECT 22.3000 53.5000 22.7000 53.6000 ;
	    RECT 23.1000 53.5000 23.4000 53.9000 ;
	    RECT 23.8000 56.2000 24.1000 64.8000 ;
	    RECT 27.0000 64.2000 27.3000 68.8000 ;
	    RECT 27.8000 66.8000 28.2000 67.2000 ;
	    RECT 27.8000 66.2000 28.1000 66.8000 ;
	    RECT 27.8000 65.8000 28.2000 66.2000 ;
	    RECT 28.6000 65.2000 28.9000 72.8000 ;
	    RECT 31.0000 66.2000 31.3000 72.8000 ;
	    RECT 32.6000 72.2000 32.9000 72.8000 ;
	    RECT 31.8000 71.8000 32.2000 72.2000 ;
	    RECT 32.6000 71.8000 33.0000 72.2000 ;
	    RECT 31.8000 67.2000 32.1000 71.8000 ;
	    RECT 31.8000 66.8000 32.2000 67.2000 ;
	    RECT 32.6000 66.8000 33.0000 67.2000 ;
	    RECT 33.4000 66.8000 33.8000 67.2000 ;
	    RECT 31.0000 65.8000 31.4000 66.2000 ;
	    RECT 32.6000 65.2000 32.9000 66.8000 ;
	    RECT 33.4000 66.2000 33.7000 66.8000 ;
	    RECT 35.8000 66.2000 36.1000 77.8000 ;
	    RECT 39.0000 76.8000 39.4000 77.2000 ;
	    RECT 40.6000 76.8000 41.0000 77.2000 ;
	    RECT 39.0000 76.2000 39.3000 76.8000 ;
	    RECT 40.6000 76.2000 40.9000 76.8000 ;
	    RECT 39.0000 75.8000 39.4000 76.2000 ;
	    RECT 40.6000 75.8000 41.0000 76.2000 ;
	    RECT 46.2000 76.1000 46.6000 76.2000 ;
	    RECT 47.0000 76.1000 47.4000 76.2000 ;
	    RECT 46.2000 75.8000 47.4000 76.1000 ;
	    RECT 49.4000 75.8000 49.8000 76.2000 ;
	    RECT 38.2000 74.8000 38.6000 75.2000 ;
	    RECT 42.2000 75.1000 42.6000 75.2000 ;
	    RECT 43.0000 75.1000 43.4000 75.2000 ;
	    RECT 42.2000 74.8000 43.4000 75.1000 ;
	    RECT 36.6000 74.1000 37.0000 74.2000 ;
	    RECT 37.4000 74.1000 37.8000 74.2000 ;
	    RECT 36.6000 73.8000 37.8000 74.1000 ;
	    RECT 36.6000 73.1000 37.0000 73.2000 ;
	    RECT 37.4000 73.1000 37.8000 73.2000 ;
	    RECT 36.6000 72.8000 37.8000 73.1000 ;
	    RECT 38.2000 72.2000 38.5000 74.8000 ;
	    RECT 39.8000 74.1000 40.2000 74.2000 ;
	    RECT 40.6000 74.1000 41.0000 74.2000 ;
	    RECT 39.8000 73.8000 41.0000 74.1000 ;
	    RECT 43.0000 73.8000 43.4000 74.2000 ;
	    RECT 45.4000 74.1000 45.8000 74.2000 ;
	    RECT 46.2000 74.1000 46.6000 74.2000 ;
	    RECT 45.4000 73.8000 46.6000 74.1000 ;
	    RECT 39.8000 73.1000 40.2000 73.2000 ;
	    RECT 39.8000 72.8000 40.9000 73.1000 ;
	    RECT 38.2000 71.8000 38.6000 72.2000 ;
	    RECT 38.2000 67.2000 38.5000 71.8000 ;
	    RECT 40.6000 69.2000 40.9000 72.8000 ;
	    RECT 40.6000 68.8000 41.0000 69.2000 ;
	    RECT 43.0000 68.2000 43.3000 73.8000 ;
	    RECT 49.4000 73.2000 49.7000 75.8000 ;
	    RECT 51.0000 75.2000 51.3000 77.8000 ;
	    RECT 51.0000 75.1000 51.4000 75.2000 ;
	    RECT 51.8000 75.1000 52.2000 75.2000 ;
	    RECT 51.0000 74.8000 52.2000 75.1000 ;
	    RECT 50.2000 74.1000 50.6000 74.2000 ;
	    RECT 51.0000 74.1000 51.4000 74.2000 ;
	    RECT 50.2000 73.8000 51.4000 74.1000 ;
	    RECT 51.8000 73.8000 52.2000 74.2000 ;
	    RECT 44.6000 73.1000 45.0000 73.2000 ;
	    RECT 45.4000 73.1000 45.8000 73.2000 ;
	    RECT 44.6000 72.8000 45.8000 73.1000 ;
	    RECT 49.4000 72.8000 49.8000 73.2000 ;
	    RECT 45.4000 68.2000 45.7000 72.8000 ;
	    RECT 51.8000 72.2000 52.1000 73.8000 ;
	    RECT 54.2000 73.2000 54.5000 85.8000 ;
	    RECT 56.6000 85.2000 56.9000 86.8000 ;
	    RECT 57.4000 86.2000 57.7000 86.8000 ;
	    RECT 57.4000 85.8000 57.8000 86.2000 ;
	    RECT 58.2000 86.1000 58.6000 86.2000 ;
	    RECT 59.0000 86.1000 59.4000 86.2000 ;
	    RECT 58.2000 85.8000 59.4000 86.1000 ;
	    RECT 56.6000 84.8000 57.0000 85.2000 ;
	    RECT 58.2000 84.8000 58.6000 85.2000 ;
	    RECT 59.0000 84.8000 59.4000 85.2000 ;
	    RECT 57.4000 77.8000 57.8000 78.2000 ;
	    RECT 56.6000 74.8000 57.0000 75.2000 ;
	    RECT 56.6000 74.2000 56.9000 74.8000 ;
	    RECT 57.4000 74.2000 57.7000 77.8000 ;
	    RECT 55.0000 74.1000 55.4000 74.2000 ;
	    RECT 55.8000 74.1000 56.2000 74.2000 ;
	    RECT 55.0000 73.8000 56.2000 74.1000 ;
	    RECT 56.6000 73.8000 57.0000 74.2000 ;
	    RECT 57.4000 73.8000 57.8000 74.2000 ;
	    RECT 54.2000 72.8000 54.6000 73.2000 ;
	    RECT 47.8000 72.1000 48.2000 72.2000 ;
	    RECT 48.6000 72.1000 49.0000 72.2000 ;
	    RECT 47.8000 71.8000 49.0000 72.1000 ;
	    RECT 51.8000 71.8000 52.2000 72.2000 ;
	    RECT 55.0000 71.8000 55.4000 72.2000 ;
	    RECT 54.2000 69.8000 54.6000 70.2000 ;
	    RECT 54.2000 69.2000 54.5000 69.8000 ;
	    RECT 55.0000 69.2000 55.3000 71.8000 ;
	    RECT 54.2000 68.8000 54.6000 69.2000 ;
	    RECT 55.0000 68.8000 55.4000 69.2000 ;
	    RECT 39.8000 67.8000 40.2000 68.2000 ;
	    RECT 43.0000 67.8000 43.4000 68.2000 ;
	    RECT 45.4000 67.8000 45.8000 68.2000 ;
	    RECT 54.2000 67.8000 54.6000 68.2000 ;
	    RECT 55.0000 67.8000 55.4000 68.2000 ;
	    RECT 39.8000 67.2000 40.1000 67.8000 ;
	    RECT 54.2000 67.2000 54.5000 67.8000 ;
	    RECT 37.4000 66.8000 37.8000 67.2000 ;
	    RECT 38.2000 66.8000 38.6000 67.2000 ;
	    RECT 39.8000 66.8000 40.2000 67.2000 ;
	    RECT 41.4000 67.1000 41.8000 67.2000 ;
	    RECT 42.2000 67.1000 42.6000 67.2000 ;
	    RECT 41.4000 66.8000 42.6000 67.1000 ;
	    RECT 43.0000 66.8000 43.4000 67.2000 ;
	    RECT 47.0000 66.8000 47.4000 67.2000 ;
	    RECT 54.2000 66.8000 54.6000 67.2000 ;
	    RECT 37.4000 66.2000 37.7000 66.8000 ;
	    RECT 33.4000 65.8000 33.8000 66.2000 ;
	    RECT 35.8000 65.8000 36.2000 66.2000 ;
	    RECT 37.4000 65.8000 37.8000 66.2000 ;
	    RECT 40.6000 65.8000 41.0000 66.2000 ;
	    RECT 35.8000 65.2000 36.1000 65.8000 ;
	    RECT 40.6000 65.2000 40.9000 65.8000 ;
	    RECT 43.0000 65.2000 43.3000 66.8000 ;
	    RECT 28.6000 64.8000 29.0000 65.2000 ;
	    RECT 32.6000 64.8000 33.0000 65.2000 ;
	    RECT 35.0000 64.8000 35.4000 65.2000 ;
	    RECT 35.8000 64.8000 36.2000 65.2000 ;
	    RECT 37.4000 65.1000 37.8000 65.2000 ;
	    RECT 38.2000 65.1000 38.6000 65.2000 ;
	    RECT 37.4000 64.8000 38.6000 65.1000 ;
	    RECT 40.6000 64.8000 41.0000 65.2000 ;
	    RECT 43.0000 64.8000 43.4000 65.2000 ;
	    RECT 35.0000 64.2000 35.3000 64.8000 ;
	    RECT 27.0000 63.8000 27.4000 64.2000 ;
	    RECT 33.4000 64.1000 33.8000 64.2000 ;
	    RECT 34.2000 64.1000 34.6000 64.2000 ;
	    RECT 33.4000 63.8000 34.6000 64.1000 ;
	    RECT 35.0000 63.8000 35.4000 64.2000 ;
	    RECT 31.0000 61.8000 31.4000 62.2000 ;
	    RECT 39.0000 61.8000 39.4000 62.2000 ;
	    RECT 31.0000 59.2000 31.3000 61.8000 ;
	    RECT 31.0000 58.8000 31.4000 59.2000 ;
	    RECT 33.4000 58.1000 33.8000 58.2000 ;
	    RECT 34.2000 58.1000 34.6000 58.2000 ;
	    RECT 23.8000 55.8000 24.2000 56.2000 ;
	    RECT 23.8000 54.2000 24.1000 55.8000 ;
	    RECT 23.8000 53.8000 24.2000 54.2000 ;
	    RECT 19.9000 53.2000 22.7000 53.5000 ;
	    RECT 19.9000 53.1000 20.3000 53.2000 ;
	    RECT 23.0000 53.1000 23.4000 53.5000 ;
	    RECT 24.6000 53.1000 25.0000 55.9000 ;
	    RECT 25.4000 53.8000 25.8000 54.2000 ;
	    RECT 25.4000 53.2000 25.7000 53.8000 ;
	    RECT 25.4000 52.8000 25.8000 53.2000 ;
	    RECT 23.0000 51.8000 23.4000 52.2000 ;
	    RECT 26.2000 52.1000 26.6000 57.9000 ;
	    RECT 27.0000 54.7000 27.4000 55.1000 ;
	    RECT 27.0000 52.2000 27.3000 54.7000 ;
	    RECT 27.0000 51.8000 27.4000 52.2000 ;
	    RECT 30.2000 51.8000 30.6000 52.2000 ;
	    RECT 31.0000 52.1000 31.4000 57.9000 ;
	    RECT 33.4000 57.8000 34.6000 58.1000 ;
	    RECT 39.0000 55.2000 39.3000 61.8000 ;
	    RECT 39.8000 58.8000 40.2000 59.2000 ;
	    RECT 39.8000 56.2000 40.1000 58.8000 ;
	    RECT 39.8000 55.8000 40.2000 56.2000 ;
	    RECT 34.2000 55.1000 34.6000 55.2000 ;
	    RECT 35.0000 55.1000 35.4000 55.2000 ;
	    RECT 34.2000 54.8000 35.4000 55.1000 ;
	    RECT 36.6000 54.8000 37.0000 55.2000 ;
	    RECT 39.0000 54.8000 39.4000 55.2000 ;
	    RECT 18.2000 49.8000 18.6000 50.2000 ;
	    RECT 17.4000 47.8000 17.8000 48.2000 ;
	    RECT 17.4000 47.2000 17.7000 47.8000 ;
	    RECT 15.8000 46.8000 16.2000 47.2000 ;
	    RECT 17.4000 46.8000 17.8000 47.2000 ;
	    RECT 10.2000 45.8000 10.6000 46.2000 ;
	    RECT 11.8000 45.8000 12.2000 46.2000 ;
	    RECT 12.6000 45.8000 13.0000 46.2000 ;
	    RECT 12.6000 45.2000 12.9000 45.8000 ;
	    RECT 12.6000 44.8000 13.0000 45.2000 ;
	    RECT 9.4000 35.8000 9.8000 36.2000 ;
	    RECT 9.4000 35.1000 9.7000 35.8000 ;
	    RECT 9.4000 34.7000 9.8000 35.1000 ;
	    RECT 6.2000 33.8000 6.6000 34.2000 ;
	    RECT 8.6000 33.8000 9.0000 34.2000 ;
	    RECT 6.2000 33.2000 6.5000 33.8000 ;
	    RECT 6.2000 32.8000 6.6000 33.2000 ;
	    RECT 0.6000 29.8000 1.0000 30.2000 ;
	    RECT 0.6000 29.2000 0.9000 29.8000 ;
	    RECT 0.6000 28.8000 1.0000 29.2000 ;
	    RECT 3.0000 23.1000 3.4000 28.9000 ;
	    RECT 7.0000 26.8000 7.4000 27.2000 ;
	    RECT 7.0000 26.3000 7.3000 26.8000 ;
	    RECT 7.0000 25.9000 7.4000 26.3000 ;
	    RECT 7.0000 25.8000 7.3000 25.9000 ;
	    RECT 7.8000 23.1000 8.2000 28.9000 ;
	    RECT 8.6000 27.2000 8.9000 33.8000 ;
	    RECT 10.2000 32.1000 10.6000 37.9000 ;
	    RECT 13.4000 37.8000 13.8000 38.2000 ;
	    RECT 11.8000 33.1000 12.2000 35.9000 ;
	    RECT 12.6000 33.8000 13.0000 34.2000 ;
	    RECT 12.6000 33.2000 12.9000 33.8000 ;
	    RECT 12.6000 32.8000 13.0000 33.2000 ;
	    RECT 8.6000 26.8000 9.0000 27.2000 ;
	    RECT 0.6000 12.1000 1.0000 12.2000 ;
	    RECT 1.4000 12.1000 1.8000 12.2000 ;
	    RECT 0.6000 11.8000 1.8000 12.1000 ;
	    RECT 2.2000 11.8000 2.6000 12.2000 ;
	    RECT 3.0000 12.1000 3.4000 17.9000 ;
	    RECT 6.2000 12.8000 6.6000 13.2000 ;
	    RECT 2.2000 6.2000 2.5000 11.8000 ;
	    RECT 6.2000 9.2000 6.5000 12.8000 ;
	    RECT 7.8000 12.1000 8.2000 17.9000 ;
	    RECT 8.6000 15.2000 8.9000 26.8000 ;
	    RECT 9.4000 25.1000 9.8000 27.9000 ;
	    RECT 10.2000 25.8000 10.6000 26.2000 ;
	    RECT 11.8000 25.8000 12.2000 26.2000 ;
	    RECT 10.2000 25.2000 10.5000 25.8000 ;
	    RECT 11.8000 25.2000 12.1000 25.8000 ;
	    RECT 13.4000 25.2000 13.7000 37.8000 ;
	    RECT 15.8000 35.2000 16.1000 46.8000 ;
	    RECT 16.6000 45.8000 17.0000 46.2000 ;
	    RECT 16.6000 45.2000 16.9000 45.8000 ;
	    RECT 16.6000 44.8000 17.0000 45.2000 ;
	    RECT 18.2000 36.2000 18.5000 49.8000 ;
	    RECT 20.6000 46.8000 21.0000 47.2000 ;
	    RECT 20.6000 46.2000 20.9000 46.8000 ;
	    RECT 20.6000 45.8000 21.0000 46.2000 ;
	    RECT 20.6000 45.2000 20.9000 45.8000 ;
	    RECT 20.6000 44.8000 21.0000 45.2000 ;
	    RECT 19.0000 43.8000 19.4000 44.2000 ;
	    RECT 19.0000 36.2000 19.3000 43.8000 ;
	    RECT 23.0000 39.2000 23.3000 51.8000 ;
	    RECT 25.4000 49.8000 25.8000 50.2000 ;
	    RECT 25.4000 48.2000 25.7000 49.8000 ;
	    RECT 24.6000 47.8000 25.0000 48.2000 ;
	    RECT 25.4000 47.8000 25.8000 48.2000 ;
	    RECT 28.6000 47.8000 29.0000 48.2000 ;
	    RECT 24.6000 47.2000 24.9000 47.8000 ;
	    RECT 24.6000 46.8000 25.0000 47.2000 ;
	    RECT 25.4000 46.8000 25.8000 47.2000 ;
	    RECT 23.8000 41.8000 24.2000 42.2000 ;
	    RECT 23.0000 38.8000 23.4000 39.2000 ;
	    RECT 23.8000 38.2000 24.1000 41.8000 ;
	    RECT 23.8000 37.8000 24.2000 38.2000 ;
	    RECT 22.2000 37.1000 22.6000 37.2000 ;
	    RECT 23.0000 37.1000 23.4000 37.2000 ;
	    RECT 22.2000 36.8000 23.4000 37.1000 ;
	    RECT 18.2000 35.8000 18.6000 36.2000 ;
	    RECT 19.0000 35.8000 19.4000 36.2000 ;
	    RECT 23.8000 35.8000 24.2000 36.2000 ;
	    RECT 14.2000 34.8000 14.6000 35.2000 ;
	    RECT 15.8000 34.8000 16.2000 35.2000 ;
	    RECT 19.8000 34.8000 20.2000 35.2000 ;
	    RECT 22.2000 35.1000 22.6000 35.2000 ;
	    RECT 23.0000 35.1000 23.4000 35.2000 ;
	    RECT 22.2000 34.8000 23.4000 35.1000 ;
	    RECT 14.2000 34.2000 14.5000 34.8000 ;
	    RECT 14.2000 33.8000 14.6000 34.2000 ;
	    RECT 16.6000 34.1000 17.0000 34.2000 ;
	    RECT 17.4000 34.1000 17.8000 34.2000 ;
	    RECT 16.6000 33.8000 17.8000 34.1000 ;
	    RECT 16.6000 27.2000 16.9000 33.8000 ;
	    RECT 17.4000 31.8000 17.8000 32.2000 ;
	    RECT 19.0000 31.8000 19.4000 32.2000 ;
	    RECT 16.6000 26.8000 17.0000 27.2000 ;
	    RECT 10.2000 24.8000 10.6000 25.2000 ;
	    RECT 11.8000 24.8000 12.2000 25.2000 ;
	    RECT 13.4000 24.8000 13.8000 25.2000 ;
	    RECT 11.8000 21.8000 12.2000 22.2000 ;
	    RECT 10.2000 19.1000 10.6000 19.2000 ;
	    RECT 11.0000 19.1000 11.4000 19.2000 ;
	    RECT 10.2000 18.8000 11.4000 19.1000 ;
	    RECT 11.0000 16.8000 11.4000 17.2000 ;
	    RECT 8.6000 14.8000 9.0000 15.2000 ;
	    RECT 8.6000 14.2000 8.9000 14.8000 ;
	    RECT 8.6000 13.8000 9.0000 14.2000 ;
	    RECT 9.4000 13.1000 9.8000 15.9000 ;
	    RECT 9.4000 10.8000 9.8000 11.2000 ;
	    RECT 6.2000 8.8000 6.6000 9.2000 ;
	    RECT 7.0000 8.8000 7.4000 9.2000 ;
	    RECT 7.0000 8.2000 7.3000 8.8000 ;
	    RECT 7.0000 7.8000 7.4000 8.2000 ;
	    RECT 7.8000 8.1000 8.2000 8.2000 ;
	    RECT 8.6000 8.1000 9.0000 8.2000 ;
	    RECT 7.8000 7.8000 9.0000 8.1000 ;
	    RECT 3.8000 7.1000 4.2000 7.2000 ;
	    RECT 4.6000 7.1000 5.0000 7.2000 ;
	    RECT 3.8000 6.8000 5.0000 7.1000 ;
	    RECT 5.4000 6.8000 5.8000 7.2000 ;
	    RECT 7.8000 6.8000 8.2000 7.2000 ;
	    RECT 5.4000 6.2000 5.7000 6.8000 ;
	    RECT 7.8000 6.2000 8.1000 6.8000 ;
	    RECT 9.4000 6.2000 9.7000 10.8000 ;
	    RECT 10.2000 7.8000 10.6000 8.2000 ;
	    RECT 10.2000 7.2000 10.5000 7.8000 ;
	    RECT 10.2000 6.8000 10.6000 7.2000 ;
	    RECT 2.2000 5.8000 2.6000 6.2000 ;
	    RECT 5.4000 5.8000 5.8000 6.2000 ;
	    RECT 7.8000 5.8000 8.2000 6.2000 ;
	    RECT 9.4000 5.8000 9.8000 6.2000 ;
	    RECT 11.0000 6.1000 11.3000 16.8000 ;
	    RECT 11.8000 9.2000 12.1000 21.8000 ;
	    RECT 12.6000 12.1000 13.0000 17.9000 ;
	    RECT 13.4000 17.2000 13.7000 24.8000 ;
	    RECT 16.6000 19.2000 16.9000 26.8000 ;
	    RECT 17.4000 26.2000 17.7000 31.8000 ;
	    RECT 17.4000 25.8000 17.8000 26.2000 ;
	    RECT 19.0000 25.2000 19.3000 31.8000 ;
	    RECT 19.8000 29.2000 20.1000 34.8000 ;
	    RECT 20.6000 34.1000 21.0000 34.2000 ;
	    RECT 21.4000 34.1000 21.8000 34.2000 ;
	    RECT 20.6000 33.8000 21.8000 34.1000 ;
	    RECT 19.8000 28.8000 20.2000 29.2000 ;
	    RECT 20.6000 28.8000 21.0000 29.2000 ;
	    RECT 20.6000 28.2000 20.9000 28.8000 ;
	    RECT 19.8000 27.8000 20.2000 28.2000 ;
	    RECT 20.6000 27.8000 21.0000 28.2000 ;
	    RECT 19.8000 26.2000 20.1000 27.8000 ;
	    RECT 23.8000 27.2000 24.1000 35.8000 ;
	    RECT 24.6000 30.2000 24.9000 46.8000 ;
	    RECT 25.4000 46.2000 25.7000 46.8000 ;
	    RECT 28.6000 46.2000 28.9000 47.8000 ;
	    RECT 30.2000 47.2000 30.5000 51.8000 ;
	    RECT 31.0000 49.8000 31.4000 50.2000 ;
	    RECT 30.2000 46.8000 30.6000 47.2000 ;
	    RECT 25.4000 45.8000 25.8000 46.2000 ;
	    RECT 28.6000 45.8000 29.0000 46.2000 ;
	    RECT 30.2000 45.2000 30.5000 46.8000 ;
	    RECT 31.0000 46.2000 31.3000 49.8000 ;
	    RECT 34.2000 47.2000 34.5000 54.8000 ;
	    RECT 36.6000 54.2000 36.9000 54.8000 ;
	    RECT 36.6000 53.8000 37.0000 54.2000 ;
	    RECT 36.6000 50.8000 37.0000 51.2000 ;
	    RECT 36.6000 49.2000 36.9000 50.8000 ;
	    RECT 39.0000 50.1000 39.3000 54.8000 ;
	    RECT 40.6000 54.2000 40.9000 64.8000 ;
	    RECT 47.0000 64.2000 47.3000 66.8000 ;
	    RECT 55.0000 66.2000 55.3000 67.8000 ;
	    RECT 55.8000 66.8000 56.2000 67.2000 ;
	    RECT 48.6000 65.8000 49.0000 66.2000 ;
	    RECT 53.4000 65.8000 53.8000 66.2000 ;
	    RECT 55.0000 65.8000 55.4000 66.2000 ;
	    RECT 48.6000 65.2000 48.9000 65.8000 ;
	    RECT 48.6000 64.8000 49.0000 65.2000 ;
	    RECT 53.4000 64.2000 53.7000 65.8000 ;
	    RECT 55.8000 64.2000 56.1000 66.8000 ;
	    RECT 56.6000 65.8000 57.0000 66.2000 ;
	    RECT 47.0000 63.8000 47.4000 64.2000 ;
	    RECT 53.4000 63.8000 53.8000 64.2000 ;
	    RECT 55.8000 63.8000 56.2000 64.2000 ;
	    RECT 43.8000 61.8000 44.2000 62.2000 ;
	    RECT 41.4000 55.8000 41.8000 56.2000 ;
	    RECT 43.0000 55.9000 43.4000 56.3000 ;
	    RECT 41.4000 54.2000 41.7000 55.8000 ;
	    RECT 42.2000 54.8000 42.6000 55.2000 ;
	    RECT 42.2000 54.2000 42.5000 54.8000 ;
	    RECT 43.0000 54.2000 43.3000 55.9000 ;
	    RECT 43.8000 55.2000 44.1000 61.8000 ;
	    RECT 56.6000 61.1000 56.9000 65.8000 ;
	    RECT 57.4000 65.2000 57.7000 73.8000 ;
	    RECT 57.4000 64.8000 57.8000 65.2000 ;
	    RECT 56.6000 60.8000 57.7000 61.1000 ;
	    RECT 54.2000 57.8000 54.6000 58.2000 ;
	    RECT 46.3000 55.9000 46.7000 56.3000 ;
	    RECT 43.8000 54.8000 44.2000 55.2000 ;
	    RECT 45.0000 54.2000 45.4000 54.3000 ;
	    RECT 40.6000 53.8000 41.0000 54.2000 ;
	    RECT 41.4000 53.8000 41.8000 54.2000 ;
	    RECT 42.2000 53.8000 42.6000 54.2000 ;
	    RECT 43.0000 53.9000 45.4000 54.2000 ;
	    RECT 39.8000 53.1000 40.2000 53.2000 ;
	    RECT 40.6000 53.1000 41.0000 53.2000 ;
	    RECT 39.8000 52.8000 41.0000 53.1000 ;
	    RECT 42.2000 51.2000 42.5000 53.8000 ;
	    RECT 43.0000 53.5000 43.3000 53.9000 ;
	    RECT 43.7000 53.5000 44.1000 53.6000 ;
	    RECT 45.4000 53.5000 45.8000 53.6000 ;
	    RECT 46.4000 53.5000 46.7000 55.9000 ;
	    RECT 50.1000 55.9000 50.5000 56.3000 ;
	    RECT 53.4000 55.9000 53.8000 56.3000 ;
	    RECT 47.0000 54.8000 47.4000 55.2000 ;
	    RECT 47.0000 54.2000 47.3000 54.8000 ;
	    RECT 47.0000 53.8000 47.4000 54.2000 ;
	    RECT 49.4000 53.8000 49.8000 54.2000 ;
	    RECT 43.0000 53.1000 43.4000 53.5000 ;
	    RECT 43.7000 53.2000 45.8000 53.5000 ;
	    RECT 46.3000 53.1000 46.7000 53.5000 ;
	    RECT 49.4000 53.2000 49.7000 53.8000 ;
	    RECT 50.1000 53.5000 50.4000 55.9000 ;
	    RECT 51.4000 54.2000 51.8000 54.3000 ;
	    RECT 53.5000 54.2000 53.8000 55.9000 ;
	    RECT 54.2000 55.2000 54.5000 57.8000 ;
	    RECT 54.2000 55.1000 54.6000 55.2000 ;
	    RECT 55.0000 55.1000 55.4000 55.2000 ;
	    RECT 54.2000 54.8000 55.4000 55.1000 ;
	    RECT 51.4000 53.9000 53.8000 54.2000 ;
	    RECT 51.0000 53.5000 51.4000 53.6000 ;
	    RECT 52.7000 53.5000 53.1000 53.6000 ;
	    RECT 53.5000 53.5000 53.8000 53.9000 ;
	    RECT 54.2000 54.1000 54.6000 54.2000 ;
	    RECT 54.2000 53.8000 55.3000 54.1000 ;
	    RECT 49.4000 52.8000 49.8000 53.2000 ;
	    RECT 50.1000 53.1000 50.5000 53.5000 ;
	    RECT 51.0000 53.2000 53.1000 53.5000 ;
	    RECT 53.4000 53.1000 53.8000 53.5000 ;
	    RECT 44.6000 51.8000 45.0000 52.2000 ;
	    RECT 51.0000 51.8000 51.4000 52.2000 ;
	    RECT 42.2000 50.8000 42.6000 51.2000 ;
	    RECT 39.0000 49.8000 40.1000 50.1000 ;
	    RECT 36.6000 48.8000 37.0000 49.2000 ;
	    RECT 34.2000 46.8000 34.6000 47.2000 ;
	    RECT 31.0000 45.8000 31.4000 46.2000 ;
	    RECT 33.4000 46.1000 33.8000 46.2000 ;
	    RECT 34.2000 46.1000 34.6000 46.2000 ;
	    RECT 33.4000 45.8000 34.6000 46.1000 ;
	    RECT 27.8000 44.8000 28.2000 45.2000 ;
	    RECT 30.2000 44.8000 30.6000 45.2000 ;
	    RECT 27.8000 44.2000 28.1000 44.8000 ;
	    RECT 25.4000 44.1000 25.8000 44.2000 ;
	    RECT 26.2000 44.1000 26.6000 44.2000 ;
	    RECT 25.4000 43.8000 26.6000 44.1000 ;
	    RECT 27.8000 43.8000 28.2000 44.2000 ;
	    RECT 28.6000 41.8000 29.0000 42.2000 ;
	    RECT 25.4000 36.8000 25.8000 37.2000 ;
	    RECT 25.4000 36.2000 25.7000 36.8000 ;
	    RECT 25.4000 35.8000 25.8000 36.2000 ;
	    RECT 27.8000 35.8000 28.2000 36.2000 ;
	    RECT 27.8000 35.2000 28.1000 35.8000 ;
	    RECT 28.6000 35.2000 28.9000 41.8000 ;
	    RECT 27.8000 34.8000 28.2000 35.2000 ;
	    RECT 28.6000 34.8000 29.0000 35.2000 ;
	    RECT 29.4000 34.8000 29.8000 35.2000 ;
	    RECT 28.6000 33.8000 29.0000 34.2000 ;
	    RECT 28.6000 33.2000 28.9000 33.8000 ;
	    RECT 28.6000 32.8000 29.0000 33.2000 ;
	    RECT 24.6000 29.8000 25.0000 30.2000 ;
	    RECT 26.2000 29.1000 26.6000 29.2000 ;
	    RECT 27.0000 29.1000 27.4000 29.2000 ;
	    RECT 26.2000 28.8000 27.4000 29.1000 ;
	    RECT 27.0000 27.8000 27.4000 28.2000 ;
	    RECT 20.6000 26.8000 21.0000 27.2000 ;
	    RECT 22.2000 26.8000 22.6000 27.2000 ;
	    RECT 23.8000 26.8000 24.2000 27.2000 ;
	    RECT 20.6000 26.2000 20.9000 26.8000 ;
	    RECT 19.8000 25.8000 20.2000 26.2000 ;
	    RECT 20.6000 25.8000 21.0000 26.2000 ;
	    RECT 19.0000 24.8000 19.4000 25.2000 ;
	    RECT 16.6000 18.8000 17.0000 19.2000 ;
	    RECT 13.4000 16.8000 13.8000 17.2000 ;
	    RECT 13.4000 15.8000 13.8000 16.2000 ;
	    RECT 16.6000 15.8000 17.0000 16.2000 ;
	    RECT 13.4000 15.2000 13.7000 15.8000 ;
	    RECT 13.4000 14.8000 13.8000 15.2000 ;
	    RECT 16.6000 15.1000 16.9000 15.8000 ;
	    RECT 16.6000 14.7000 17.0000 15.1000 ;
	    RECT 16.6000 11.8000 17.0000 12.2000 ;
	    RECT 17.4000 12.1000 17.8000 17.9000 ;
	    RECT 19.0000 17.1000 19.3000 24.8000 ;
	    RECT 22.2000 21.1000 22.5000 26.8000 ;
	    RECT 25.4000 25.8000 25.8000 26.2000 ;
	    RECT 24.6000 24.8000 25.0000 25.2000 ;
	    RECT 24.6000 24.2000 24.9000 24.8000 ;
	    RECT 24.6000 23.8000 25.0000 24.2000 ;
	    RECT 22.2000 20.8000 23.3000 21.1000 ;
	    RECT 23.0000 19.2000 23.3000 20.8000 ;
	    RECT 25.4000 19.2000 25.7000 25.8000 ;
	    RECT 27.0000 22.2000 27.3000 27.8000 ;
	    RECT 27.0000 21.8000 27.4000 22.2000 ;
	    RECT 28.6000 21.8000 29.0000 22.2000 ;
	    RECT 23.0000 18.8000 23.4000 19.2000 ;
	    RECT 25.4000 18.8000 25.8000 19.2000 ;
	    RECT 27.8000 18.8000 28.2000 19.2000 ;
	    RECT 18.2000 16.8000 19.3000 17.1000 ;
	    RECT 20.6000 17.8000 21.0000 18.2000 ;
	    RECT 20.6000 17.2000 20.9000 17.8000 ;
	    RECT 20.6000 16.8000 21.0000 17.2000 ;
	    RECT 25.4000 16.8000 25.8000 17.2000 ;
	    RECT 26.2000 16.8000 26.6000 17.2000 ;
	    RECT 16.6000 9.2000 16.9000 11.8000 ;
	    RECT 18.2000 11.2000 18.5000 16.8000 ;
	    RECT 19.0000 13.1000 19.4000 15.9000 ;
	    RECT 19.8000 15.8000 20.2000 16.2000 ;
	    RECT 22.2000 15.8000 22.6000 16.2000 ;
	    RECT 19.8000 15.2000 20.1000 15.8000 ;
	    RECT 22.2000 15.2000 22.5000 15.8000 ;
	    RECT 25.4000 15.2000 25.7000 16.8000 ;
	    RECT 26.2000 16.2000 26.5000 16.8000 ;
	    RECT 26.2000 15.8000 26.6000 16.2000 ;
	    RECT 19.8000 14.8000 20.2000 15.2000 ;
	    RECT 21.4000 14.8000 21.8000 15.2000 ;
	    RECT 22.2000 14.8000 22.6000 15.2000 ;
	    RECT 25.4000 14.8000 25.8000 15.2000 ;
	    RECT 21.4000 13.2000 21.7000 14.8000 ;
	    RECT 21.4000 12.8000 21.8000 13.2000 ;
	    RECT 23.8000 12.8000 24.2000 13.2000 ;
	    RECT 23.8000 11.2000 24.1000 12.8000 ;
	    RECT 18.2000 10.8000 18.6000 11.2000 ;
	    RECT 23.8000 10.8000 24.2000 11.2000 ;
	    RECT 18.2000 10.2000 18.5000 10.8000 ;
	    RECT 18.2000 9.8000 18.6000 10.2000 ;
	    RECT 23.8000 9.8000 24.2000 10.2000 ;
	    RECT 11.8000 8.8000 12.2000 9.2000 ;
	    RECT 15.8000 8.8000 16.2000 9.2000 ;
	    RECT 16.6000 8.8000 17.0000 9.2000 ;
	    RECT 15.8000 8.2000 16.1000 8.8000 ;
	    RECT 15.8000 8.1000 16.2000 8.2000 ;
	    RECT 16.6000 8.1000 17.0000 8.2000 ;
	    RECT 15.8000 7.8000 17.0000 8.1000 ;
	    RECT 18.2000 7.2000 18.5000 9.8000 ;
	    RECT 22.2000 8.8000 22.6000 9.2000 ;
	    RECT 22.2000 8.2000 22.5000 8.8000 ;
	    RECT 22.2000 7.8000 22.6000 8.2000 ;
	    RECT 11.8000 7.1000 12.2000 7.2000 ;
	    RECT 12.6000 7.1000 13.0000 7.2000 ;
	    RECT 11.8000 6.8000 13.0000 7.1000 ;
	    RECT 18.2000 6.8000 18.6000 7.2000 ;
	    RECT 23.0000 6.8000 23.4000 7.2000 ;
	    RECT 23.0000 6.2000 23.3000 6.8000 ;
	    RECT 23.8000 6.2000 24.1000 9.8000 ;
	    RECT 10.2000 5.8000 11.3000 6.1000 ;
	    RECT 15.8000 5.8000 16.2000 6.2000 ;
	    RECT 18.2000 6.1000 18.6000 6.2000 ;
	    RECT 19.0000 6.1000 19.4000 6.2000 ;
	    RECT 18.2000 5.8000 19.4000 6.1000 ;
	    RECT 23.0000 5.8000 23.4000 6.2000 ;
	    RECT 23.8000 5.8000 24.2000 6.2000 ;
	    RECT 10.2000 5.2000 10.5000 5.8000 ;
	    RECT 15.8000 5.2000 16.1000 5.8000 ;
	    RECT 25.4000 5.2000 25.7000 14.8000 ;
	    RECT 27.8000 13.2000 28.1000 18.8000 ;
	    RECT 28.6000 18.2000 28.9000 21.8000 ;
	    RECT 28.6000 17.8000 29.0000 18.2000 ;
	    RECT 28.6000 15.8000 29.0000 16.2000 ;
	    RECT 28.6000 15.2000 28.9000 15.8000 ;
	    RECT 29.4000 15.2000 29.7000 34.8000 ;
	    RECT 30.2000 34.2000 30.5000 44.8000 ;
	    RECT 31.0000 35.2000 31.3000 45.8000 ;
	    RECT 34.2000 44.8000 34.6000 45.2000 ;
	    RECT 34.2000 44.2000 34.5000 44.8000 ;
	    RECT 34.2000 43.8000 34.6000 44.2000 ;
	    RECT 39.0000 43.1000 39.4000 48.9000 ;
	    RECT 35.8000 41.8000 36.2000 42.2000 ;
	    RECT 35.8000 39.2000 36.1000 41.8000 ;
	    RECT 35.8000 38.8000 36.2000 39.2000 ;
	    RECT 34.2000 37.8000 34.6000 38.2000 ;
	    RECT 32.6000 35.8000 33.0000 36.2000 ;
	    RECT 32.6000 35.2000 32.9000 35.8000 ;
	    RECT 34.2000 35.2000 34.5000 37.8000 ;
	    RECT 39.8000 37.1000 40.1000 49.8000 ;
	    RECT 43.0000 45.9000 43.4000 46.3000 ;
	    RECT 43.0000 45.2000 43.3000 45.9000 ;
	    RECT 43.0000 44.8000 43.4000 45.2000 ;
	    RECT 43.8000 43.1000 44.2000 48.9000 ;
	    RECT 44.6000 46.2000 44.9000 51.8000 ;
	    RECT 44.6000 45.8000 45.0000 46.2000 ;
	    RECT 45.4000 45.1000 45.8000 47.9000 ;
	    RECT 47.8000 45.1000 48.2000 47.9000 ;
	    RECT 49.4000 43.1000 49.8000 48.9000 ;
	    RECT 51.0000 46.2000 51.3000 51.8000 ;
	    RECT 51.0000 45.8000 51.4000 46.2000 ;
	    RECT 53.4000 45.8000 53.8000 46.2000 ;
	    RECT 53.4000 42.2000 53.7000 45.8000 ;
	    RECT 54.2000 43.1000 54.6000 48.9000 ;
	    RECT 55.0000 48.2000 55.3000 53.8000 ;
	    RECT 56.6000 51.8000 57.0000 52.2000 ;
	    RECT 55.0000 47.8000 55.4000 48.2000 ;
	    RECT 56.6000 45.2000 56.9000 51.8000 ;
	    RECT 57.4000 46.2000 57.7000 60.8000 ;
	    RECT 58.2000 57.2000 58.5000 84.8000 ;
	    RECT 59.0000 84.2000 59.3000 84.8000 ;
	    RECT 59.0000 83.8000 59.4000 84.2000 ;
	    RECT 59.0000 70.2000 59.3000 83.8000 ;
	    RECT 59.8000 77.2000 60.1000 87.8000 ;
	    RECT 66.2000 87.2000 66.5000 113.8000 ;
	    RECT 67.8000 113.2000 68.1000 113.8000 ;
	    RECT 67.8000 112.8000 68.2000 113.2000 ;
	    RECT 68.6000 109.2000 68.9000 114.8000 ;
	    RECT 71.0000 113.1000 71.4000 115.9000 ;
	    RECT 72.6000 112.1000 73.0000 117.9000 ;
	    RECT 73.4000 115.8000 73.8000 116.2000 ;
	    RECT 73.4000 115.1000 73.7000 115.8000 ;
	    RECT 73.4000 114.7000 73.8000 115.1000 ;
	    RECT 75.0000 113.8000 75.4000 114.2000 ;
	    RECT 75.0000 111.2000 75.3000 113.8000 ;
	    RECT 77.4000 112.1000 77.8000 117.9000 ;
	    RECT 95.9000 115.9000 96.3000 116.3000 ;
	    RECT 99.0000 115.9000 99.4000 116.3000 ;
	    RECT 83.0000 114.8000 83.4000 115.2000 ;
	    RECT 85.4000 114.8000 85.8000 115.2000 ;
	    RECT 87.0000 115.1000 87.4000 115.2000 ;
	    RECT 87.8000 115.1000 88.2000 115.2000 ;
	    RECT 87.0000 114.8000 88.2000 115.1000 ;
	    RECT 89.4000 115.1000 89.8000 115.2000 ;
	    RECT 90.2000 115.1000 90.6000 115.2000 ;
	    RECT 89.4000 114.8000 90.6000 115.1000 ;
	    RECT 92.6000 114.8000 93.0000 115.2000 ;
	    RECT 78.2000 114.1000 78.6000 114.2000 ;
	    RECT 79.0000 114.1000 79.4000 114.2000 ;
	    RECT 78.2000 113.8000 79.4000 114.1000 ;
	    RECT 75.0000 110.8000 75.4000 111.2000 ;
	    RECT 78.2000 110.8000 78.6000 111.2000 ;
	    RECT 67.8000 108.8000 68.2000 109.2000 ;
	    RECT 68.6000 108.8000 69.0000 109.2000 ;
	    RECT 74.2000 108.8000 74.6000 109.2000 ;
	    RECT 67.0000 107.8000 67.4000 108.2000 ;
	    RECT 67.0000 107.2000 67.3000 107.8000 ;
	    RECT 67.0000 106.8000 67.4000 107.2000 ;
	    RECT 67.0000 105.8000 67.4000 106.2000 ;
	    RECT 67.0000 105.2000 67.3000 105.8000 ;
	    RECT 67.0000 104.8000 67.4000 105.2000 ;
	    RECT 67.8000 95.2000 68.1000 108.8000 ;
	    RECT 74.2000 108.2000 74.5000 108.8000 ;
	    RECT 68.5000 107.5000 68.9000 107.9000 ;
	    RECT 69.4000 107.5000 71.5000 107.8000 ;
	    RECT 71.8000 107.5000 72.2000 107.9000 ;
	    RECT 68.5000 105.1000 68.8000 107.5000 ;
	    RECT 69.4000 107.4000 69.8000 107.5000 ;
	    RECT 71.1000 107.4000 71.5000 107.5000 ;
	    RECT 71.9000 107.1000 72.2000 107.5000 ;
	    RECT 69.8000 106.8000 72.2000 107.1000 ;
	    RECT 69.8000 106.7000 70.2000 106.8000 ;
	    RECT 71.9000 105.1000 72.2000 106.8000 ;
	    RECT 74.2000 107.8000 74.6000 108.2000 ;
	    RECT 68.5000 104.7000 68.9000 105.1000 ;
	    RECT 71.8000 104.7000 72.2000 105.1000 ;
	    RECT 72.6000 105.8000 73.0000 106.2000 ;
	    RECT 72.6000 105.2000 72.9000 105.8000 ;
	    RECT 72.6000 104.8000 73.0000 105.2000 ;
	    RECT 74.2000 104.2000 74.5000 107.8000 ;
	    RECT 74.2000 103.8000 74.6000 104.2000 ;
	    RECT 77.4000 103.1000 77.8000 108.9000 ;
	    RECT 78.2000 106.2000 78.5000 110.8000 ;
	    RECT 78.2000 105.8000 78.6000 106.2000 ;
	    RECT 79.8000 106.1000 80.2000 106.2000 ;
	    RECT 80.6000 106.1000 81.0000 106.2000 ;
	    RECT 79.8000 105.8000 81.0000 106.1000 ;
	    RECT 68.6000 99.8000 69.0000 100.2000 ;
	    RECT 67.8000 94.8000 68.2000 95.2000 ;
	    RECT 67.8000 93.8000 68.2000 94.2000 ;
	    RECT 63.8000 87.1000 64.2000 87.2000 ;
	    RECT 64.6000 87.1000 65.0000 87.2000 ;
	    RECT 63.8000 86.8000 65.0000 87.1000 ;
	    RECT 65.4000 86.8000 65.8000 87.2000 ;
	    RECT 66.2000 86.8000 66.6000 87.2000 ;
	    RECT 65.4000 86.2000 65.7000 86.8000 ;
	    RECT 60.6000 85.8000 61.0000 86.2000 ;
	    RECT 63.0000 86.1000 63.4000 86.2000 ;
	    RECT 63.0000 85.8000 64.1000 86.1000 ;
	    RECT 60.6000 85.2000 60.9000 85.8000 ;
	    RECT 63.8000 85.2000 64.1000 85.8000 ;
	    RECT 65.4000 85.8000 65.8000 86.2000 ;
	    RECT 65.4000 85.2000 65.7000 85.8000 ;
	    RECT 60.6000 84.8000 61.0000 85.2000 ;
	    RECT 63.8000 84.8000 64.2000 85.2000 ;
	    RECT 65.4000 84.8000 65.8000 85.2000 ;
	    RECT 61.4000 79.1000 61.8000 79.2000 ;
	    RECT 62.2000 79.1000 62.6000 79.2000 ;
	    RECT 61.4000 78.8000 62.6000 79.1000 ;
	    RECT 59.8000 76.8000 60.2000 77.2000 ;
	    RECT 63.8000 72.1000 64.2000 77.9000 ;
	    RECT 66.2000 75.2000 66.5000 86.8000 ;
	    RECT 67.8000 78.2000 68.1000 93.8000 ;
	    RECT 68.6000 93.2000 68.9000 99.8000 ;
	    RECT 70.2000 95.1000 70.6000 95.2000 ;
	    RECT 71.0000 95.1000 71.4000 95.2000 ;
	    RECT 70.2000 94.8000 71.4000 95.1000 ;
	    RECT 71.8000 94.8000 72.2000 95.2000 ;
	    RECT 68.6000 92.8000 69.0000 93.2000 ;
	    RECT 70.2000 92.8000 70.6000 93.2000 ;
	    RECT 70.2000 89.2000 70.5000 92.8000 ;
	    RECT 71.8000 90.2000 72.1000 94.8000 ;
	    RECT 72.6000 93.1000 73.0000 95.9000 ;
	    RECT 74.2000 92.1000 74.6000 97.9000 ;
	    RECT 75.0000 95.8000 75.4000 96.2000 ;
	    RECT 75.0000 95.1000 75.3000 95.8000 ;
	    RECT 78.2000 95.2000 78.5000 105.8000 ;
	    RECT 82.2000 103.1000 82.6000 108.9000 ;
	    RECT 81.4000 99.8000 81.8000 100.2000 ;
	    RECT 81.4000 99.2000 81.7000 99.8000 ;
	    RECT 81.4000 98.8000 81.8000 99.2000 ;
	    RECT 75.0000 94.7000 75.4000 95.1000 ;
	    RECT 78.2000 94.8000 78.6000 95.2000 ;
	    RECT 71.8000 89.8000 72.2000 90.2000 ;
	    RECT 70.2000 88.8000 70.6000 89.2000 ;
	    RECT 75.0000 89.1000 75.4000 89.2000 ;
	    RECT 75.8000 89.1000 76.2000 89.2000 ;
	    RECT 75.0000 88.8000 76.2000 89.1000 ;
	    RECT 78.2000 88.2000 78.5000 94.8000 ;
	    RECT 79.0000 92.1000 79.4000 97.9000 ;
	    RECT 82.2000 94.8000 82.6000 95.2000 ;
	    RECT 82.2000 94.2000 82.5000 94.8000 ;
	    RECT 82.2000 93.8000 82.6000 94.2000 ;
	    RECT 73.3000 87.5000 73.7000 87.9000 ;
	    RECT 74.2000 87.5000 76.3000 87.8000 ;
	    RECT 76.6000 87.5000 77.0000 87.9000 ;
	    RECT 69.4000 86.8000 69.8000 87.2000 ;
	    RECT 71.8000 87.1000 72.2000 87.2000 ;
	    RECT 72.6000 87.1000 73.0000 87.2000 ;
	    RECT 71.8000 86.8000 73.0000 87.1000 ;
	    RECT 69.4000 86.2000 69.7000 86.8000 ;
	    RECT 69.4000 85.8000 69.8000 86.2000 ;
	    RECT 71.8000 85.8000 72.2000 86.2000 ;
	    RECT 68.6000 84.8000 69.0000 85.2000 ;
	    RECT 68.6000 84.2000 68.9000 84.8000 ;
	    RECT 68.6000 83.8000 69.0000 84.2000 ;
	    RECT 71.8000 81.2000 72.1000 85.8000 ;
	    RECT 73.3000 85.1000 73.6000 87.5000 ;
	    RECT 74.2000 87.4000 74.6000 87.5000 ;
	    RECT 75.9000 87.4000 76.3000 87.5000 ;
	    RECT 76.7000 87.1000 77.0000 87.5000 ;
	    RECT 74.6000 86.8000 77.0000 87.1000 ;
	    RECT 77.4000 87.8000 77.8000 88.2000 ;
	    RECT 78.2000 87.8000 78.6000 88.2000 ;
	    RECT 77.4000 87.2000 77.7000 87.8000 ;
	    RECT 77.4000 87.1000 77.8000 87.2000 ;
	    RECT 77.4000 86.8000 78.5000 87.1000 ;
	    RECT 74.6000 86.7000 75.0000 86.8000 ;
	    RECT 74.2000 85.8000 74.6000 86.2000 ;
	    RECT 73.3000 84.7000 73.7000 85.1000 ;
	    RECT 71.8000 80.8000 72.2000 81.2000 ;
	    RECT 74.2000 79.2000 74.5000 85.8000 ;
	    RECT 76.7000 85.1000 77.0000 86.8000 ;
	    RECT 76.6000 84.7000 77.0000 85.1000 ;
	    RECT 78.2000 84.2000 78.5000 86.8000 ;
	    RECT 78.2000 83.8000 78.6000 84.2000 ;
	    RECT 79.8000 83.8000 80.2000 84.2000 ;
	    RECT 74.2000 78.8000 74.6000 79.2000 ;
	    RECT 67.8000 77.8000 68.2000 78.2000 ;
	    RECT 66.2000 74.8000 66.6000 75.2000 ;
	    RECT 67.8000 74.7000 68.2000 75.1000 ;
	    RECT 59.0000 69.8000 59.4000 70.2000 ;
	    RECT 67.8000 69.2000 68.1000 74.7000 ;
	    RECT 68.6000 72.1000 69.0000 77.9000 ;
	    RECT 77.4000 77.8000 77.8000 78.2000 ;
	    RECT 79.0000 77.8000 79.4000 78.2000 ;
	    RECT 69.4000 75.8000 69.8000 76.2000 ;
	    RECT 71.8000 75.9000 72.2000 76.3000 ;
	    RECT 75.1000 75.9000 75.5000 76.3000 ;
	    RECT 69.4000 74.2000 69.7000 75.8000 ;
	    RECT 69.4000 73.8000 69.8000 74.2000 ;
	    RECT 70.2000 73.1000 70.6000 75.9000 ;
	    RECT 71.8000 74.2000 72.1000 75.9000 ;
	    RECT 73.8000 74.2000 74.2000 74.3000 ;
	    RECT 71.0000 73.8000 71.4000 74.2000 ;
	    RECT 71.8000 73.9000 74.2000 74.2000 ;
	    RECT 71.0000 72.2000 71.3000 73.8000 ;
	    RECT 71.8000 73.5000 72.1000 73.9000 ;
	    RECT 72.5000 73.5000 72.9000 73.6000 ;
	    RECT 74.2000 73.5000 74.6000 73.6000 ;
	    RECT 75.2000 73.5000 75.5000 75.9000 ;
	    RECT 71.8000 73.1000 72.2000 73.5000 ;
	    RECT 72.5000 73.2000 74.6000 73.5000 ;
	    RECT 75.1000 73.1000 75.5000 73.5000 ;
	    RECT 76.6000 74.8000 77.0000 75.2000 ;
	    RECT 71.0000 71.8000 71.4000 72.2000 ;
	    RECT 72.6000 71.8000 73.0000 72.2000 ;
	    RECT 72.6000 71.2000 72.9000 71.8000 ;
	    RECT 72.6000 70.8000 73.0000 71.2000 ;
	    RECT 72.6000 69.2000 72.9000 70.8000 ;
	    RECT 76.6000 70.2000 76.9000 74.8000 ;
	    RECT 76.6000 69.8000 77.0000 70.2000 ;
	    RECT 60.6000 68.8000 61.0000 69.2000 ;
	    RECT 67.8000 68.8000 68.2000 69.2000 ;
	    RECT 72.6000 68.8000 73.0000 69.2000 ;
	    RECT 59.0000 65.1000 59.4000 65.2000 ;
	    RECT 59.8000 65.1000 60.2000 65.2000 ;
	    RECT 59.0000 64.8000 60.2000 65.1000 ;
	    RECT 60.6000 65.1000 60.9000 68.8000 ;
	    RECT 66.1000 67.5000 66.5000 67.9000 ;
	    RECT 67.0000 67.5000 69.1000 67.8000 ;
	    RECT 69.4000 67.5000 69.8000 67.9000 ;
	    RECT 61.4000 67.1000 61.8000 67.2000 ;
	    RECT 62.2000 67.1000 62.6000 67.2000 ;
	    RECT 61.4000 66.8000 62.6000 67.1000 ;
	    RECT 64.6000 67.1000 65.0000 67.2000 ;
	    RECT 65.4000 67.1000 65.8000 67.2000 ;
	    RECT 64.6000 66.8000 65.8000 67.1000 ;
	    RECT 64.6000 65.8000 65.0000 66.2000 ;
	    RECT 61.4000 65.1000 61.8000 65.2000 ;
	    RECT 60.6000 64.8000 61.8000 65.1000 ;
	    RECT 63.0000 64.8000 63.4000 65.2000 ;
	    RECT 63.0000 64.2000 63.3000 64.8000 ;
	    RECT 63.0000 63.8000 63.4000 64.2000 ;
	    RECT 58.2000 56.8000 58.6000 57.2000 ;
	    RECT 58.2000 56.2000 58.5000 56.8000 ;
	    RECT 58.2000 55.8000 58.6000 56.2000 ;
	    RECT 64.6000 55.2000 64.9000 65.8000 ;
	    RECT 66.1000 65.1000 66.4000 67.5000 ;
	    RECT 67.0000 67.4000 67.4000 67.5000 ;
	    RECT 68.7000 67.4000 69.1000 67.5000 ;
	    RECT 69.5000 67.1000 69.8000 67.5000 ;
	    RECT 67.4000 66.8000 69.8000 67.1000 ;
	    RECT 70.2000 67.8000 70.6000 68.2000 ;
	    RECT 70.2000 67.2000 70.5000 67.8000 ;
	    RECT 70.2000 66.8000 70.6000 67.2000 ;
	    RECT 67.4000 66.7000 67.8000 66.8000 ;
	    RECT 69.5000 65.1000 69.8000 66.8000 ;
	    RECT 77.4000 66.2000 77.7000 77.8000 ;
	    RECT 79.0000 74.2000 79.3000 77.8000 ;
	    RECT 79.8000 76.2000 80.1000 83.8000 ;
	    RECT 80.6000 83.1000 81.0000 88.9000 ;
	    RECT 82.2000 85.2000 82.5000 93.8000 ;
	    RECT 82.2000 84.8000 82.6000 85.2000 ;
	    RECT 83.0000 79.2000 83.3000 114.8000 ;
	    RECT 83.8000 105.1000 84.2000 107.9000 ;
	    RECT 84.6000 105.8000 85.0000 106.2000 ;
	    RECT 84.6000 100.2000 84.9000 105.8000 ;
	    RECT 84.6000 99.8000 85.0000 100.2000 ;
	    RECT 85.4000 94.2000 85.7000 114.8000 ;
	    RECT 87.8000 110.8000 88.2000 111.2000 ;
	    RECT 87.0000 105.1000 87.4000 107.9000 ;
	    RECT 87.8000 107.2000 88.1000 110.8000 ;
	    RECT 92.6000 109.2000 92.9000 114.8000 ;
	    RECT 95.0000 114.1000 95.4000 114.2000 ;
	    RECT 94.2000 113.8000 95.4000 114.1000 ;
	    RECT 87.8000 106.8000 88.2000 107.2000 ;
	    RECT 88.6000 103.1000 89.0000 108.9000 ;
	    RECT 92.6000 108.8000 93.0000 109.2000 ;
	    RECT 92.6000 107.8000 93.0000 108.2000 ;
	    RECT 92.6000 107.2000 92.9000 107.8000 ;
	    RECT 92.6000 106.8000 93.0000 107.2000 ;
	    RECT 89.4000 105.9000 89.8000 106.3000 ;
	    RECT 89.4000 99.2000 89.7000 105.9000 ;
	    RECT 93.4000 103.1000 93.8000 108.9000 ;
	    RECT 94.2000 108.1000 94.5000 113.8000 ;
	    RECT 95.9000 113.5000 96.2000 115.9000 ;
	    RECT 96.5000 114.9000 96.9000 115.3000 ;
	    RECT 96.6000 114.2000 96.9000 114.9000 ;
	    RECT 99.1000 114.2000 99.4000 115.9000 ;
	    RECT 96.6000 113.9000 99.4000 114.2000 ;
	    RECT 96.6000 113.5000 97.0000 113.6000 ;
	    RECT 98.3000 113.5000 98.7000 113.6000 ;
	    RECT 99.1000 113.5000 99.4000 113.9000 ;
	    RECT 95.9000 113.2000 98.7000 113.5000 ;
	    RECT 95.9000 113.1000 96.3000 113.2000 ;
	    RECT 99.0000 113.1000 99.4000 113.5000 ;
	    RECT 102.2000 114.8000 102.6000 115.2000 ;
	    RECT 104.6000 114.8000 105.0000 115.2000 ;
	    RECT 97.4000 112.1000 97.8000 112.2000 ;
	    RECT 98.2000 112.1000 98.6000 112.2000 ;
	    RECT 97.4000 111.8000 98.6000 112.1000 ;
	    RECT 101.4000 111.8000 101.8000 112.2000 ;
	    RECT 95.0000 109.1000 95.4000 109.2000 ;
	    RECT 95.8000 109.1000 96.2000 109.2000 ;
	    RECT 95.0000 108.8000 96.2000 109.1000 ;
	    RECT 94.2000 107.8000 95.3000 108.1000 ;
	    RECT 95.0000 99.2000 95.3000 107.8000 ;
	    RECT 96.6000 104.8000 97.0000 105.2000 ;
	    RECT 98.2000 105.1000 98.6000 107.9000 ;
	    RECT 99.0000 106.8000 99.4000 107.2000 ;
	    RECT 99.0000 106.2000 99.3000 106.8000 ;
	    RECT 99.0000 105.8000 99.4000 106.2000 ;
	    RECT 96.6000 99.2000 96.9000 104.8000 ;
	    RECT 99.8000 103.1000 100.2000 108.9000 ;
	    RECT 101.4000 106.2000 101.7000 111.8000 ;
	    RECT 102.2000 110.2000 102.5000 114.8000 ;
	    RECT 104.6000 111.2000 104.9000 114.8000 ;
	    RECT 107.0000 114.1000 107.4000 114.2000 ;
	    RECT 107.8000 114.1000 108.2000 114.2000 ;
	    RECT 107.0000 113.8000 108.2000 114.1000 ;
	    RECT 109.4000 113.8000 109.8000 114.2000 ;
	    RECT 108.6000 111.8000 109.0000 112.2000 ;
	    RECT 108.6000 111.2000 108.9000 111.8000 ;
	    RECT 104.6000 110.8000 105.0000 111.2000 ;
	    RECT 106.2000 110.8000 106.6000 111.2000 ;
	    RECT 108.6000 110.8000 109.0000 111.2000 ;
	    RECT 102.2000 109.8000 102.6000 110.2000 ;
	    RECT 101.4000 105.8000 101.8000 106.2000 ;
	    RECT 104.6000 103.1000 105.0000 108.9000 ;
	    RECT 105.4000 106.8000 105.8000 107.2000 ;
	    RECT 89.4000 98.8000 89.8000 99.2000 ;
	    RECT 95.0000 98.8000 95.4000 99.2000 ;
	    RECT 96.6000 98.8000 97.0000 99.2000 ;
	    RECT 90.2000 96.8000 90.6000 97.2000 ;
	    RECT 90.2000 95.2000 90.5000 96.8000 ;
	    RECT 91.0000 95.8000 91.4000 96.2000 ;
	    RECT 91.0000 95.2000 91.3000 95.8000 ;
	    RECT 86.2000 94.8000 86.6000 95.2000 ;
	    RECT 87.8000 94.8000 88.2000 95.2000 ;
	    RECT 90.2000 94.8000 90.6000 95.2000 ;
	    RECT 91.0000 94.8000 91.4000 95.2000 ;
	    RECT 91.8000 94.8000 92.2000 95.2000 ;
	    RECT 94.2000 94.8000 94.6000 95.2000 ;
	    RECT 86.2000 94.2000 86.5000 94.8000 ;
	    RECT 85.4000 93.8000 85.8000 94.2000 ;
	    RECT 86.2000 93.8000 86.6000 94.2000 ;
	    RECT 87.8000 89.2000 88.1000 94.8000 ;
	    RECT 91.8000 94.2000 92.1000 94.8000 ;
	    RECT 89.4000 93.8000 89.8000 94.2000 ;
	    RECT 91.8000 93.8000 92.2000 94.2000 ;
	    RECT 89.4000 89.2000 89.7000 93.8000 ;
	    RECT 94.2000 93.2000 94.5000 94.8000 ;
	    RECT 97.4000 93.8000 97.8000 94.2000 ;
	    RECT 97.4000 93.2000 97.7000 93.8000 ;
	    RECT 94.2000 92.8000 94.6000 93.2000 ;
	    RECT 97.4000 92.8000 97.8000 93.2000 ;
	    RECT 103.8000 92.8000 104.2000 93.2000 ;
	    RECT 95.0000 91.8000 95.4000 92.2000 ;
	    RECT 96.6000 91.8000 97.0000 92.2000 ;
	    RECT 83.8000 88.8000 84.2000 89.2000 ;
	    RECT 83.8000 86.2000 84.1000 88.8000 ;
	    RECT 83.8000 85.8000 84.2000 86.2000 ;
	    RECT 85.4000 83.1000 85.8000 88.9000 ;
	    RECT 87.8000 88.8000 88.2000 89.2000 ;
	    RECT 89.4000 88.8000 89.8000 89.2000 ;
	    RECT 95.0000 88.2000 95.3000 91.8000 ;
	    RECT 96.6000 89.2000 96.9000 91.8000 ;
	    RECT 103.0000 90.8000 103.4000 91.2000 ;
	    RECT 103.0000 89.2000 103.3000 90.8000 ;
	    RECT 96.6000 88.8000 97.0000 89.2000 ;
	    RECT 103.0000 88.8000 103.4000 89.2000 ;
	    RECT 86.2000 87.8000 86.6000 88.2000 ;
	    RECT 86.2000 87.2000 86.5000 87.8000 ;
	    RECT 86.2000 86.8000 86.6000 87.2000 ;
	    RECT 87.0000 85.1000 87.4000 87.9000 ;
	    RECT 95.0000 87.8000 95.4000 88.2000 ;
	    RECT 103.8000 87.2000 104.1000 92.8000 ;
	    RECT 104.6000 92.1000 105.0000 97.9000 ;
	    RECT 105.4000 95.2000 105.7000 106.8000 ;
	    RECT 105.4000 94.8000 105.8000 95.2000 ;
	    RECT 105.4000 91.2000 105.7000 94.8000 ;
	    RECT 105.4000 90.8000 105.8000 91.2000 ;
	    RECT 95.0000 87.1000 95.4000 87.2000 ;
	    RECT 95.8000 87.1000 96.2000 87.2000 ;
	    RECT 95.0000 86.8000 96.2000 87.1000 ;
	    RECT 99.0000 86.8000 99.4000 87.2000 ;
	    RECT 103.8000 86.8000 104.2000 87.2000 ;
	    RECT 87.8000 85.8000 88.2000 86.2000 ;
	    RECT 98.2000 85.8000 98.6000 86.2000 ;
	    RECT 87.0000 82.8000 87.4000 83.2000 ;
	    RECT 87.0000 79.2000 87.3000 82.8000 ;
	    RECT 87.8000 81.2000 88.1000 85.8000 ;
	    RECT 98.2000 85.2000 98.5000 85.8000 ;
	    RECT 95.8000 84.8000 96.2000 85.2000 ;
	    RECT 96.6000 84.8000 97.0000 85.2000 ;
	    RECT 98.2000 84.8000 98.6000 85.2000 ;
	    RECT 93.4000 83.8000 93.8000 84.2000 ;
	    RECT 87.8000 80.8000 88.2000 81.2000 ;
	    RECT 93.4000 79.2000 93.7000 83.8000 ;
	    RECT 83.0000 78.8000 83.4000 79.2000 ;
	    RECT 87.0000 78.8000 87.4000 79.2000 ;
	    RECT 93.4000 78.8000 93.8000 79.2000 ;
	    RECT 83.0000 77.8000 83.4000 78.2000 ;
	    RECT 89.4000 77.8000 89.8000 78.2000 ;
	    RECT 81.4000 76.8000 81.8000 77.2000 ;
	    RECT 81.4000 76.2000 81.7000 76.8000 ;
	    RECT 79.8000 75.8000 80.2000 76.2000 ;
	    RECT 80.6000 75.8000 81.0000 76.2000 ;
	    RECT 81.4000 75.8000 81.8000 76.2000 ;
	    RECT 79.0000 73.8000 79.4000 74.2000 ;
	    RECT 78.2000 73.1000 78.6000 73.2000 ;
	    RECT 79.0000 73.1000 79.4000 73.2000 ;
	    RECT 78.2000 72.8000 79.4000 73.1000 ;
	    RECT 79.8000 71.8000 80.2000 72.2000 ;
	    RECT 78.2000 68.8000 78.6000 69.2000 ;
	    RECT 66.1000 64.7000 66.5000 65.1000 ;
	    RECT 69.4000 64.7000 69.8000 65.1000 ;
	    RECT 70.2000 65.8000 70.6000 66.2000 ;
	    RECT 77.4000 65.8000 77.8000 66.2000 ;
	    RECT 70.2000 55.2000 70.5000 65.8000 ;
	    RECT 77.4000 65.2000 77.7000 65.8000 ;
	    RECT 77.4000 64.8000 77.8000 65.2000 ;
	    RECT 78.2000 62.2000 78.5000 68.8000 ;
	    RECT 79.0000 67.8000 79.4000 68.2000 ;
	    RECT 79.0000 67.2000 79.3000 67.8000 ;
	    RECT 79.0000 66.8000 79.4000 67.2000 ;
	    RECT 78.2000 61.8000 78.6000 62.2000 ;
	    RECT 78.2000 60.8000 78.6000 61.2000 ;
	    RECT 72.6000 55.8000 73.0000 56.2000 ;
	    RECT 63.0000 54.8000 63.4000 55.2000 ;
	    RECT 64.6000 54.8000 65.0000 55.2000 ;
	    RECT 69.4000 55.1000 69.8000 55.2000 ;
	    RECT 70.2000 55.1000 70.6000 55.2000 ;
	    RECT 69.4000 54.8000 70.6000 55.1000 ;
	    RECT 71.0000 54.8000 71.4000 55.2000 ;
	    RECT 59.8000 54.1000 60.2000 54.4000 ;
	    RECT 60.6000 54.1000 61.0000 54.2000 ;
	    RECT 59.8000 53.8000 61.0000 54.1000 ;
	    RECT 61.4000 52.8000 61.8000 53.2000 ;
	    RECT 61.4000 48.2000 61.7000 52.8000 ;
	    RECT 63.0000 52.2000 63.3000 54.8000 ;
	    RECT 71.0000 54.2000 71.3000 54.8000 ;
	    RECT 63.8000 54.1000 64.2000 54.2000 ;
	    RECT 64.6000 54.1000 65.0000 54.2000 ;
	    RECT 63.8000 53.8000 65.0000 54.1000 ;
	    RECT 67.0000 53.8000 67.4000 54.2000 ;
	    RECT 67.8000 54.1000 68.2000 54.2000 ;
	    RECT 68.6000 54.1000 69.0000 54.2000 ;
	    RECT 67.8000 53.8000 69.0000 54.1000 ;
	    RECT 70.2000 54.1000 70.6000 54.2000 ;
	    RECT 71.0000 54.1000 71.4000 54.2000 ;
	    RECT 70.2000 53.8000 71.4000 54.1000 ;
	    RECT 64.6000 52.8000 65.0000 53.2000 ;
	    RECT 65.4000 53.1000 65.8000 53.2000 ;
	    RECT 66.2000 53.1000 66.6000 53.2000 ;
	    RECT 65.4000 52.8000 66.6000 53.1000 ;
	    RECT 63.0000 51.8000 63.4000 52.2000 ;
	    RECT 64.6000 50.2000 64.9000 52.8000 ;
	    RECT 64.6000 49.8000 65.0000 50.2000 ;
	    RECT 67.0000 48.2000 67.3000 53.8000 ;
	    RECT 61.4000 47.8000 61.8000 48.2000 ;
	    RECT 62.2000 48.1000 62.6000 48.2000 ;
	    RECT 63.0000 48.1000 63.4000 48.2000 ;
	    RECT 62.2000 47.8000 63.4000 48.1000 ;
	    RECT 65.4000 47.8000 65.8000 48.2000 ;
	    RECT 66.2000 48.1000 66.6000 48.2000 ;
	    RECT 67.0000 48.1000 67.4000 48.2000 ;
	    RECT 66.2000 47.8000 67.4000 48.1000 ;
	    RECT 63.8000 47.1000 64.2000 47.2000 ;
	    RECT 64.6000 47.1000 65.0000 47.2000 ;
	    RECT 63.8000 46.8000 65.0000 47.1000 ;
	    RECT 57.4000 45.8000 57.8000 46.2000 ;
	    RECT 59.8000 45.8000 60.2000 46.2000 ;
	    RECT 56.6000 44.8000 57.0000 45.2000 ;
	    RECT 59.8000 44.2000 60.1000 45.8000 ;
	    RECT 63.8000 44.8000 64.2000 45.2000 ;
	    RECT 56.6000 44.1000 57.0000 44.2000 ;
	    RECT 57.4000 44.1000 57.8000 44.2000 ;
	    RECT 56.6000 43.8000 57.8000 44.1000 ;
	    RECT 59.8000 43.8000 60.2000 44.2000 ;
	    RECT 53.4000 41.8000 53.8000 42.2000 ;
	    RECT 52.6000 38.8000 53.0000 39.2000 ;
	    RECT 55.0000 38.8000 55.4000 39.2000 ;
	    RECT 39.0000 36.8000 40.1000 37.1000 ;
	    RECT 40.6000 36.8000 41.0000 37.2000 ;
	    RECT 39.0000 36.2000 39.3000 36.8000 ;
	    RECT 40.6000 36.2000 40.9000 36.8000 ;
	    RECT 52.6000 36.2000 52.9000 38.8000 ;
	    RECT 37.4000 35.8000 37.8000 36.2000 ;
	    RECT 38.8000 35.8000 39.3000 36.2000 ;
	    RECT 39.8000 35.8000 40.2000 36.2000 ;
	    RECT 40.6000 35.8000 41.0000 36.2000 ;
	    RECT 45.4000 35.8000 45.8000 36.2000 ;
	    RECT 46.2000 35.8000 46.6000 36.2000 ;
	    RECT 51.8000 35.8000 52.2000 36.2000 ;
	    RECT 52.6000 35.8000 53.0000 36.2000 ;
	    RECT 37.4000 35.2000 37.7000 35.8000 ;
	    RECT 39.8000 35.2000 40.1000 35.8000 ;
	    RECT 31.0000 34.8000 31.4000 35.2000 ;
	    RECT 32.6000 34.8000 33.0000 35.2000 ;
	    RECT 33.4000 35.1000 33.8000 35.2000 ;
	    RECT 34.2000 35.1000 34.6000 35.2000 ;
	    RECT 33.4000 34.8000 34.6000 35.1000 ;
	    RECT 37.4000 34.8000 37.8000 35.2000 ;
	    RECT 39.8000 34.8000 40.2000 35.2000 ;
	    RECT 30.2000 33.8000 30.6000 34.2000 ;
	    RECT 37.4000 33.8000 37.8000 34.2000 ;
	    RECT 42.2000 33.8000 42.6000 34.2000 ;
	    RECT 31.0000 32.8000 31.4000 33.2000 ;
	    RECT 32.6000 33.1000 33.0000 33.2000 ;
	    RECT 33.4000 33.1000 33.8000 33.2000 ;
	    RECT 32.6000 32.8000 33.8000 33.1000 ;
	    RECT 31.0000 31.2000 31.3000 32.8000 ;
	    RECT 35.8000 31.8000 36.2000 32.2000 ;
	    RECT 31.0000 30.8000 31.4000 31.2000 ;
	    RECT 31.8000 29.8000 32.2000 30.2000 ;
	    RECT 31.8000 27.2000 32.1000 29.8000 ;
	    RECT 35.8000 29.1000 36.1000 31.8000 ;
	    RECT 37.4000 31.2000 37.7000 33.8000 ;
	    RECT 42.2000 32.2000 42.5000 33.8000 ;
	    RECT 45.4000 33.2000 45.7000 35.8000 ;
	    RECT 46.2000 35.2000 46.5000 35.8000 ;
	    RECT 51.8000 35.2000 52.1000 35.8000 ;
	    RECT 46.2000 34.8000 46.6000 35.2000 ;
	    RECT 51.0000 34.8000 51.4000 35.2000 ;
	    RECT 51.8000 34.8000 52.2000 35.2000 ;
	    RECT 52.6000 35.1000 53.0000 35.2000 ;
	    RECT 53.4000 35.1000 53.8000 35.2000 ;
	    RECT 52.6000 34.8000 53.8000 35.1000 ;
	    RECT 43.0000 32.8000 43.4000 33.2000 ;
	    RECT 45.4000 32.8000 45.8000 33.2000 ;
	    RECT 46.2000 32.8000 46.6000 33.2000 ;
	    RECT 43.0000 32.2000 43.3000 32.8000 ;
	    RECT 42.2000 31.8000 42.6000 32.2000 ;
	    RECT 43.0000 31.8000 43.4000 32.2000 ;
	    RECT 44.6000 31.8000 45.0000 32.2000 ;
	    RECT 37.4000 30.8000 37.8000 31.2000 ;
	    RECT 35.8000 28.8000 36.9000 29.1000 ;
	    RECT 35.8000 27.8000 36.2000 28.2000 ;
	    RECT 35.8000 27.2000 36.1000 27.8000 ;
	    RECT 36.6000 27.2000 36.9000 28.8000 ;
	    RECT 31.0000 26.8000 31.4000 27.2000 ;
	    RECT 31.8000 26.8000 32.2000 27.2000 ;
	    RECT 35.8000 26.8000 36.2000 27.2000 ;
	    RECT 36.6000 26.8000 37.0000 27.2000 ;
	    RECT 31.0000 26.2000 31.3000 26.8000 ;
	    RECT 31.0000 25.8000 31.4000 26.2000 ;
	    RECT 31.8000 25.8000 32.2000 26.2000 ;
	    RECT 31.8000 25.1000 32.1000 25.8000 ;
	    RECT 31.0000 24.8000 32.1000 25.1000 ;
	    RECT 37.4000 25.1000 37.7000 30.8000 ;
	    RECT 41.4000 27.8000 41.8000 28.2000 ;
	    RECT 43.8000 27.8000 44.2000 28.2000 ;
	    RECT 41.4000 27.2000 41.7000 27.8000 ;
	    RECT 43.8000 27.2000 44.1000 27.8000 ;
	    RECT 44.6000 27.2000 44.9000 31.8000 ;
	    RECT 45.4000 28.2000 45.7000 32.8000 ;
	    RECT 46.2000 31.2000 46.5000 32.8000 ;
	    RECT 46.2000 30.8000 46.6000 31.2000 ;
	    RECT 46.2000 30.2000 46.5000 30.8000 ;
	    RECT 46.2000 29.8000 46.6000 30.2000 ;
	    RECT 51.0000 28.2000 51.3000 34.8000 ;
	    RECT 55.0000 34.2000 55.3000 38.8000 ;
	    RECT 58.2000 37.8000 58.6000 38.2000 ;
	    RECT 63.0000 37.8000 63.4000 38.2000 ;
	    RECT 58.2000 36.2000 58.5000 37.8000 ;
	    RECT 58.2000 35.8000 58.6000 36.2000 ;
	    RECT 57.4000 35.1000 57.8000 35.2000 ;
	    RECT 58.2000 35.1000 58.6000 35.2000 ;
	    RECT 57.4000 34.8000 58.6000 35.1000 ;
	    RECT 59.8000 34.8000 60.2000 35.2000 ;
	    RECT 60.6000 35.1000 61.0000 35.2000 ;
	    RECT 61.4000 35.1000 61.8000 35.2000 ;
	    RECT 60.6000 34.8000 61.8000 35.1000 ;
	    RECT 51.8000 33.8000 52.2000 34.2000 ;
	    RECT 55.0000 33.8000 55.4000 34.2000 ;
	    RECT 51.8000 33.2000 52.1000 33.8000 ;
	    RECT 57.4000 33.2000 57.7000 34.8000 ;
	    RECT 59.8000 33.2000 60.1000 34.8000 ;
	    RECT 60.6000 33.8000 61.0000 34.2000 ;
	    RECT 51.8000 32.8000 52.2000 33.2000 ;
	    RECT 57.4000 32.8000 57.8000 33.2000 ;
	    RECT 59.8000 32.8000 60.2000 33.2000 ;
	    RECT 59.8000 32.2000 60.1000 32.8000 ;
	    RECT 60.6000 32.2000 60.9000 33.8000 ;
	    RECT 58.2000 31.8000 58.6000 32.2000 ;
	    RECT 59.8000 31.8000 60.2000 32.2000 ;
	    RECT 60.6000 31.8000 61.0000 32.2000 ;
	    RECT 51.8000 29.8000 52.2000 30.2000 ;
	    RECT 45.4000 27.8000 45.8000 28.2000 ;
	    RECT 51.0000 27.8000 51.4000 28.2000 ;
	    RECT 51.8000 27.2000 52.1000 29.8000 ;
	    RECT 53.4000 28.1000 53.8000 28.2000 ;
	    RECT 54.2000 28.1000 54.6000 28.2000 ;
	    RECT 53.4000 27.8000 54.6000 28.1000 ;
	    RECT 38.2000 27.1000 38.6000 27.2000 ;
	    RECT 39.0000 27.1000 39.4000 27.2000 ;
	    RECT 38.2000 26.8000 39.4000 27.1000 ;
	    RECT 39.8000 26.8000 40.2000 27.2000 ;
	    RECT 41.4000 26.8000 41.8000 27.2000 ;
	    RECT 42.2000 26.8000 42.6000 27.2000 ;
	    RECT 43.8000 26.8000 44.2000 27.2000 ;
	    RECT 44.6000 26.8000 45.0000 27.2000 ;
	    RECT 47.8000 26.8000 48.2000 27.2000 ;
	    RECT 51.8000 26.8000 52.2000 27.2000 ;
	    RECT 53.4000 27.1000 53.8000 27.2000 ;
	    RECT 54.2000 27.1000 54.6000 27.2000 ;
	    RECT 53.4000 26.8000 54.6000 27.1000 ;
	    RECT 57.4000 26.8000 57.8000 27.2000 ;
	    RECT 39.8000 25.2000 40.1000 26.8000 ;
	    RECT 42.2000 26.2000 42.5000 26.8000 ;
	    RECT 40.6000 25.8000 41.0000 26.2000 ;
	    RECT 42.2000 25.8000 42.6000 26.2000 ;
	    RECT 44.6000 26.1000 45.0000 26.2000 ;
	    RECT 45.4000 26.1000 45.8000 26.2000 ;
	    RECT 44.6000 25.8000 45.8000 26.1000 ;
	    RECT 37.4000 24.8000 38.5000 25.1000 ;
	    RECT 39.8000 24.8000 40.2000 25.2000 ;
	    RECT 31.0000 23.2000 31.3000 24.8000 ;
	    RECT 32.6000 23.8000 33.0000 24.2000 ;
	    RECT 31.0000 22.8000 31.4000 23.2000 ;
	    RECT 31.0000 19.2000 31.3000 22.8000 ;
	    RECT 32.6000 19.2000 32.9000 23.8000 ;
	    RECT 31.0000 18.8000 31.4000 19.2000 ;
	    RECT 32.6000 18.8000 33.0000 19.2000 ;
	    RECT 30.2000 16.8000 30.6000 17.2000 ;
	    RECT 28.6000 14.8000 29.0000 15.2000 ;
	    RECT 29.4000 14.8000 29.8000 15.2000 ;
	    RECT 30.2000 14.2000 30.5000 16.8000 ;
	    RECT 32.6000 16.2000 32.9000 18.8000 ;
	    RECT 31.0000 16.1000 31.4000 16.2000 ;
	    RECT 31.8000 16.1000 32.2000 16.2000 ;
	    RECT 31.0000 15.8000 32.2000 16.1000 ;
	    RECT 32.6000 15.8000 33.0000 16.2000 ;
	    RECT 31.8000 14.8000 32.2000 15.2000 ;
	    RECT 35.0000 14.8000 35.4000 15.2000 ;
	    RECT 35.8000 14.8000 36.2000 15.2000 ;
	    RECT 37.4000 14.8000 37.8000 15.2000 ;
	    RECT 31.8000 14.2000 32.1000 14.8000 ;
	    RECT 35.0000 14.2000 35.3000 14.8000 ;
	    RECT 30.2000 13.8000 30.6000 14.2000 ;
	    RECT 31.8000 13.8000 32.2000 14.2000 ;
	    RECT 35.0000 13.8000 35.4000 14.2000 ;
	    RECT 35.8000 13.2000 36.1000 14.8000 ;
	    RECT 37.4000 14.2000 37.7000 14.8000 ;
	    RECT 37.4000 13.8000 37.8000 14.2000 ;
	    RECT 27.8000 12.8000 28.2000 13.2000 ;
	    RECT 35.8000 13.1000 36.2000 13.2000 ;
	    RECT 36.6000 13.1000 37.0000 13.2000 ;
	    RECT 35.8000 12.8000 37.0000 13.1000 ;
	    RECT 27.0000 11.8000 27.4000 12.2000 ;
	    RECT 36.6000 11.8000 37.0000 12.2000 ;
	    RECT 27.0000 9.2000 27.3000 11.8000 ;
	    RECT 36.6000 11.2000 36.9000 11.8000 ;
	    RECT 36.6000 10.8000 37.0000 11.2000 ;
	    RECT 35.0000 9.8000 35.4000 10.2000 ;
	    RECT 27.0000 8.8000 27.4000 9.2000 ;
	    RECT 29.4000 8.8000 29.8000 9.2000 ;
	    RECT 29.4000 7.2000 29.7000 8.8000 ;
	    RECT 35.0000 7.2000 35.3000 9.8000 ;
	    RECT 38.2000 9.2000 38.5000 24.8000 ;
	    RECT 39.0000 12.8000 39.4000 13.2000 ;
	    RECT 37.4000 9.1000 37.8000 9.2000 ;
	    RECT 38.2000 9.1000 38.6000 9.2000 ;
	    RECT 37.4000 8.8000 38.6000 9.1000 ;
	    RECT 27.8000 7.1000 28.2000 7.2000 ;
	    RECT 28.6000 7.1000 29.0000 7.2000 ;
	    RECT 27.8000 6.8000 29.0000 7.1000 ;
	    RECT 29.4000 6.8000 29.8000 7.2000 ;
	    RECT 35.0000 6.8000 35.4000 7.2000 ;
	    RECT 29.4000 6.1000 29.8000 6.2000 ;
	    RECT 30.2000 6.1000 30.6000 6.2000 ;
	    RECT 29.4000 5.8000 30.6000 6.1000 ;
	    RECT 32.6000 5.8000 33.0000 6.2000 ;
	    RECT 38.2000 6.1000 38.6000 6.2000 ;
	    RECT 39.0000 6.1000 39.3000 12.8000 ;
	    RECT 40.6000 11.2000 40.9000 25.8000 ;
	    RECT 47.8000 24.2000 48.1000 26.8000 ;
	    RECT 57.4000 26.2000 57.7000 26.8000 ;
	    RECT 48.6000 25.8000 49.0000 26.2000 ;
	    RECT 50.2000 25.8000 50.6000 26.2000 ;
	    RECT 51.0000 25.8000 51.4000 26.2000 ;
	    RECT 51.8000 25.8000 52.2000 26.2000 ;
	    RECT 52.6000 26.1000 53.0000 26.2000 ;
	    RECT 53.4000 26.1000 53.8000 26.2000 ;
	    RECT 52.6000 25.8000 53.8000 26.1000 ;
	    RECT 55.8000 26.1000 56.2000 26.2000 ;
	    RECT 56.6000 26.1000 57.0000 26.2000 ;
	    RECT 55.8000 25.8000 57.0000 26.1000 ;
	    RECT 57.4000 25.8000 57.8000 26.2000 ;
	    RECT 58.2000 26.1000 58.5000 31.8000 ;
	    RECT 59.8000 27.8000 60.2000 28.2000 ;
	    RECT 59.8000 27.2000 60.1000 27.8000 ;
	    RECT 59.8000 26.8000 60.2000 27.2000 ;
	    RECT 61.4000 27.1000 61.7000 34.8000 ;
	    RECT 63.0000 34.2000 63.3000 37.8000 ;
	    RECT 63.8000 34.2000 64.1000 44.8000 ;
	    RECT 65.4000 36.2000 65.7000 47.8000 ;
	    RECT 67.0000 47.1000 67.4000 47.2000 ;
	    RECT 67.8000 47.1000 68.1000 53.8000 ;
	    RECT 72.6000 52.2000 72.9000 55.8000 ;
	    RECT 75.0000 55.1000 75.4000 55.2000 ;
	    RECT 74.2000 54.8000 75.4000 55.1000 ;
	    RECT 74.2000 53.2000 74.5000 54.8000 ;
	    RECT 78.2000 54.2000 78.5000 60.8000 ;
	    RECT 75.0000 54.1000 75.4000 54.2000 ;
	    RECT 75.8000 54.1000 76.2000 54.2000 ;
	    RECT 75.0000 53.8000 76.2000 54.1000 ;
	    RECT 78.2000 53.8000 78.6000 54.2000 ;
	    RECT 74.2000 52.8000 74.6000 53.2000 ;
	    RECT 75.8000 53.1000 76.2000 53.2000 ;
	    RECT 76.6000 53.1000 77.0000 53.2000 ;
	    RECT 75.8000 52.8000 77.0000 53.1000 ;
	    RECT 77.4000 52.8000 77.8000 53.2000 ;
	    RECT 77.4000 52.2000 77.7000 52.8000 ;
	    RECT 71.8000 51.8000 72.2000 52.2000 ;
	    RECT 72.6000 51.8000 73.0000 52.2000 ;
	    RECT 74.2000 51.8000 74.6000 52.2000 ;
	    RECT 77.4000 51.8000 77.8000 52.2000 ;
	    RECT 67.0000 46.8000 68.1000 47.1000 ;
	    RECT 69.4000 49.8000 69.8000 50.2000 ;
	    RECT 69.4000 47.2000 69.7000 49.8000 ;
	    RECT 71.0000 47.8000 71.4000 48.2000 ;
	    RECT 71.0000 47.2000 71.3000 47.8000 ;
	    RECT 69.4000 46.8000 69.8000 47.2000 ;
	    RECT 71.0000 46.8000 71.4000 47.2000 ;
	    RECT 68.6000 45.8000 69.0000 46.2000 ;
	    RECT 68.6000 45.2000 68.9000 45.8000 ;
	    RECT 68.6000 44.8000 69.0000 45.2000 ;
	    RECT 67.0000 37.8000 67.4000 38.2000 ;
	    RECT 65.4000 35.8000 65.8000 36.2000 ;
	    RECT 63.0000 33.8000 63.4000 34.2000 ;
	    RECT 63.8000 33.8000 64.2000 34.2000 ;
	    RECT 65.4000 28.2000 65.7000 35.8000 ;
	    RECT 67.0000 33.2000 67.3000 37.8000 ;
	    RECT 69.4000 35.2000 69.7000 46.8000 ;
	    RECT 68.6000 34.8000 69.0000 35.2000 ;
	    RECT 69.4000 34.8000 69.8000 35.2000 ;
	    RECT 68.6000 33.2000 68.9000 34.8000 ;
	    RECT 66.2000 32.8000 66.6000 33.2000 ;
	    RECT 67.0000 32.8000 67.4000 33.2000 ;
	    RECT 67.8000 32.8000 68.2000 33.2000 ;
	    RECT 68.6000 32.8000 69.0000 33.2000 ;
	    RECT 71.0000 32.8000 71.4000 33.2000 ;
	    RECT 66.2000 32.2000 66.5000 32.8000 ;
	    RECT 67.8000 32.2000 68.1000 32.8000 ;
	    RECT 71.0000 32.2000 71.3000 32.8000 ;
	    RECT 66.2000 31.8000 66.6000 32.2000 ;
	    RECT 67.8000 31.8000 68.2000 32.2000 ;
	    RECT 69.4000 31.8000 69.8000 32.2000 ;
	    RECT 71.0000 31.8000 71.4000 32.2000 ;
	    RECT 66.2000 28.2000 66.5000 31.8000 ;
	    RECT 65.4000 27.8000 65.8000 28.2000 ;
	    RECT 66.2000 27.8000 66.6000 28.2000 ;
	    RECT 60.6000 26.8000 61.7000 27.1000 ;
	    RECT 67.8000 27.2000 68.1000 31.8000 ;
	    RECT 69.4000 31.2000 69.7000 31.8000 ;
	    RECT 69.4000 30.8000 69.8000 31.2000 ;
	    RECT 71.8000 27.2000 72.1000 51.8000 ;
	    RECT 72.6000 48.2000 72.9000 51.8000 ;
	    RECT 73.4000 48.8000 73.8000 49.2000 ;
	    RECT 73.4000 48.2000 73.7000 48.8000 ;
	    RECT 72.6000 47.8000 73.0000 48.2000 ;
	    RECT 73.4000 47.8000 73.8000 48.2000 ;
	    RECT 73.4000 46.2000 73.7000 47.8000 ;
	    RECT 73.4000 45.8000 73.8000 46.2000 ;
	    RECT 74.2000 44.2000 74.5000 51.8000 ;
	    RECT 75.0000 48.1000 75.4000 48.2000 ;
	    RECT 75.8000 48.1000 76.2000 48.2000 ;
	    RECT 75.0000 47.8000 76.2000 48.1000 ;
	    RECT 77.4000 47.8000 77.8000 48.2000 ;
	    RECT 75.0000 46.8000 75.4000 47.2000 ;
	    RECT 75.8000 46.8000 76.2000 47.2000 ;
	    RECT 75.0000 46.2000 75.3000 46.8000 ;
	    RECT 75.8000 46.2000 76.1000 46.8000 ;
	    RECT 75.0000 45.8000 75.4000 46.2000 ;
	    RECT 75.8000 45.8000 76.2000 46.2000 ;
	    RECT 77.4000 45.2000 77.7000 47.8000 ;
	    RECT 77.4000 44.8000 77.8000 45.2000 ;
	    RECT 74.2000 43.8000 74.6000 44.2000 ;
	    RECT 77.4000 39.2000 77.7000 44.8000 ;
	    RECT 75.8000 39.1000 76.2000 39.2000 ;
	    RECT 76.6000 39.1000 77.0000 39.2000 ;
	    RECT 75.8000 38.8000 77.0000 39.1000 ;
	    RECT 77.4000 38.8000 77.8000 39.2000 ;
	    RECT 72.6000 36.8000 73.0000 37.2000 ;
	    RECT 75.0000 36.8000 75.4000 37.2000 ;
	    RECT 76.6000 37.1000 77.0000 37.2000 ;
	    RECT 77.4000 37.1000 77.8000 37.2000 ;
	    RECT 76.6000 36.8000 77.8000 37.1000 ;
	    RECT 72.6000 36.2000 72.9000 36.8000 ;
	    RECT 75.0000 36.2000 75.3000 36.8000 ;
	    RECT 72.6000 35.8000 73.0000 36.2000 ;
	    RECT 75.0000 35.8000 75.4000 36.2000 ;
	    RECT 72.6000 30.2000 72.9000 35.8000 ;
	    RECT 78.2000 35.2000 78.5000 53.8000 ;
	    RECT 79.8000 52.2000 80.1000 71.8000 ;
	    RECT 80.6000 70.2000 80.9000 75.8000 ;
	    RECT 83.0000 75.2000 83.3000 77.8000 ;
	    RECT 89.4000 77.2000 89.7000 77.8000 ;
	    RECT 86.2000 76.8000 86.6000 77.2000 ;
	    RECT 88.6000 76.8000 89.0000 77.2000 ;
	    RECT 89.4000 76.8000 89.8000 77.2000 ;
	    RECT 84.6000 75.8000 85.0000 76.2000 ;
	    RECT 85.4000 75.8000 85.8000 76.2000 ;
	    RECT 84.6000 75.2000 84.9000 75.8000 ;
	    RECT 85.4000 75.2000 85.7000 75.8000 ;
	    RECT 83.0000 74.8000 83.4000 75.2000 ;
	    RECT 84.6000 74.8000 85.0000 75.2000 ;
	    RECT 85.4000 74.8000 85.8000 75.2000 ;
	    RECT 83.8000 73.8000 84.2000 74.2000 ;
	    RECT 81.4000 72.8000 81.8000 73.2000 ;
	    RECT 81.4000 72.2000 81.7000 72.8000 ;
	    RECT 81.4000 71.8000 81.8000 72.2000 ;
	    RECT 80.6000 69.8000 81.0000 70.2000 ;
	    RECT 81.4000 69.2000 81.7000 71.8000 ;
	    RECT 83.0000 69.8000 83.4000 70.2000 ;
	    RECT 83.0000 69.2000 83.3000 69.8000 ;
	    RECT 81.4000 68.8000 81.8000 69.2000 ;
	    RECT 83.0000 68.8000 83.4000 69.2000 ;
	    RECT 83.8000 68.2000 84.1000 73.8000 ;
	    RECT 84.6000 70.2000 84.9000 74.8000 ;
	    RECT 86.2000 70.2000 86.5000 76.8000 ;
	    RECT 88.6000 76.2000 88.9000 76.8000 ;
	    RECT 95.8000 76.2000 96.1000 84.8000 ;
	    RECT 96.6000 79.2000 96.9000 84.8000 ;
	    RECT 99.0000 83.2000 99.3000 86.8000 ;
	    RECT 99.0000 82.8000 99.4000 83.2000 ;
	    RECT 99.8000 82.8000 100.2000 83.2000 ;
	    RECT 99.0000 79.2000 99.3000 82.8000 ;
	    RECT 96.6000 78.8000 97.0000 79.2000 ;
	    RECT 99.0000 78.8000 99.4000 79.2000 ;
	    RECT 97.4000 77.1000 97.8000 77.2000 ;
	    RECT 98.2000 77.1000 98.6000 77.2000 ;
	    RECT 97.4000 76.8000 98.6000 77.1000 ;
	    RECT 99.0000 76.8000 99.4000 77.2000 ;
	    RECT 99.0000 76.2000 99.3000 76.8000 ;
	    RECT 88.6000 75.8000 89.0000 76.2000 ;
	    RECT 90.2000 76.1000 90.6000 76.2000 ;
	    RECT 91.0000 76.1000 91.4000 76.2000 ;
	    RECT 90.2000 75.8000 91.4000 76.1000 ;
	    RECT 95.8000 75.8000 96.2000 76.2000 ;
	    RECT 99.0000 75.8000 99.4000 76.2000 ;
	    RECT 88.6000 75.1000 89.0000 75.2000 ;
	    RECT 89.4000 75.1000 89.8000 75.2000 ;
	    RECT 88.6000 74.8000 89.8000 75.1000 ;
	    RECT 91.0000 74.8000 91.4000 75.2000 ;
	    RECT 91.8000 74.8000 92.2000 75.2000 ;
	    RECT 94.2000 74.8000 94.6000 75.2000 ;
	    RECT 96.6000 74.8000 97.0000 75.2000 ;
	    RECT 89.4000 74.2000 89.7000 74.8000 ;
	    RECT 89.4000 73.8000 89.8000 74.2000 ;
	    RECT 91.0000 71.2000 91.3000 74.8000 ;
	    RECT 91.8000 74.2000 92.1000 74.8000 ;
	    RECT 91.8000 73.8000 92.2000 74.2000 ;
	    RECT 94.2000 72.2000 94.5000 74.8000 ;
	    RECT 96.6000 73.2000 96.9000 74.8000 ;
	    RECT 96.6000 72.8000 97.0000 73.2000 ;
	    RECT 94.2000 71.8000 94.6000 72.2000 ;
	    RECT 91.0000 70.8000 91.4000 71.2000 ;
	    RECT 84.6000 69.8000 85.0000 70.2000 ;
	    RECT 86.2000 69.8000 86.6000 70.2000 ;
	    RECT 87.0000 69.1000 87.4000 69.2000 ;
	    RECT 87.8000 69.1000 88.2000 69.2000 ;
	    RECT 87.0000 68.8000 88.2000 69.1000 ;
	    RECT 91.0000 68.8000 91.4000 69.2000 ;
	    RECT 94.2000 68.8000 94.6000 69.2000 ;
	    RECT 91.0000 68.2000 91.3000 68.8000 ;
	    RECT 94.2000 68.2000 94.5000 68.8000 ;
	    RECT 82.2000 67.8000 82.6000 68.2000 ;
	    RECT 83.8000 67.8000 84.2000 68.2000 ;
	    RECT 86.2000 67.8000 86.6000 68.2000 ;
	    RECT 91.0000 67.8000 91.4000 68.2000 ;
	    RECT 94.2000 67.8000 94.6000 68.2000 ;
	    RECT 82.2000 67.2000 82.5000 67.8000 ;
	    RECT 86.2000 67.2000 86.5000 67.8000 ;
	    RECT 80.6000 66.8000 81.0000 67.2000 ;
	    RECT 82.2000 66.8000 82.6000 67.2000 ;
	    RECT 84.6000 67.1000 85.0000 67.2000 ;
	    RECT 85.4000 67.1000 85.8000 67.2000 ;
	    RECT 84.6000 66.8000 85.8000 67.1000 ;
	    RECT 86.2000 66.8000 86.6000 67.2000 ;
	    RECT 88.6000 67.1000 89.0000 67.2000 ;
	    RECT 89.4000 67.1000 89.8000 67.2000 ;
	    RECT 88.6000 66.8000 89.8000 67.1000 ;
	    RECT 92.6000 66.8000 93.0000 67.2000 ;
	    RECT 95.8000 66.8000 96.2000 67.2000 ;
	    RECT 80.6000 66.2000 80.9000 66.8000 ;
	    RECT 80.6000 66.1000 81.0000 66.2000 ;
	    RECT 81.4000 66.1000 81.8000 66.2000 ;
	    RECT 80.6000 65.8000 81.8000 66.1000 ;
	    RECT 84.6000 66.1000 85.0000 66.2000 ;
	    RECT 85.4000 66.1000 85.8000 66.2000 ;
	    RECT 84.6000 65.8000 85.8000 66.1000 ;
	    RECT 84.6000 61.8000 85.0000 62.2000 ;
	    RECT 84.6000 57.2000 84.9000 61.8000 ;
	    RECT 84.6000 56.8000 85.0000 57.2000 ;
	    RECT 84.6000 56.2000 84.9000 56.8000 ;
	    RECT 84.6000 55.8000 85.0000 56.2000 ;
	    RECT 86.2000 55.2000 86.5000 66.8000 ;
	    RECT 92.6000 66.2000 92.9000 66.8000 ;
	    RECT 95.8000 66.2000 96.1000 66.8000 ;
	    RECT 90.2000 65.8000 90.6000 66.2000 ;
	    RECT 91.0000 65.8000 91.4000 66.2000 ;
	    RECT 92.6000 65.8000 93.0000 66.2000 ;
	    RECT 95.8000 65.8000 96.2000 66.2000 ;
	    RECT 90.2000 65.2000 90.5000 65.8000 ;
	    RECT 87.0000 65.1000 87.4000 65.2000 ;
	    RECT 87.8000 65.1000 88.2000 65.2000 ;
	    RECT 87.0000 64.8000 88.2000 65.1000 ;
	    RECT 90.2000 64.8000 90.6000 65.2000 ;
	    RECT 87.8000 58.8000 88.2000 59.2000 ;
	    RECT 87.8000 58.2000 88.1000 58.8000 ;
	    RECT 87.8000 57.8000 88.2000 58.2000 ;
	    RECT 90.2000 56.2000 90.5000 64.8000 ;
	    RECT 90.2000 55.8000 90.6000 56.2000 ;
	    RECT 91.0000 55.2000 91.3000 65.8000 ;
	    RECT 96.6000 63.2000 96.9000 72.8000 ;
	    RECT 99.8000 69.2000 100.1000 82.8000 ;
	    RECT 103.8000 78.2000 104.1000 86.8000 ;
	    RECT 106.2000 82.2000 106.5000 110.8000 ;
	    RECT 109.4000 110.2000 109.7000 113.8000 ;
	    RECT 111.8000 113.1000 112.2000 115.9000 ;
	    RECT 112.6000 113.8000 113.0000 114.2000 ;
	    RECT 111.0000 111.8000 111.4000 112.2000 ;
	    RECT 107.0000 109.8000 107.4000 110.2000 ;
	    RECT 109.4000 109.8000 109.8000 110.2000 ;
	    RECT 107.0000 109.2000 107.3000 109.8000 ;
	    RECT 107.0000 108.8000 107.4000 109.2000 ;
	    RECT 107.8000 108.8000 108.2000 109.2000 ;
	    RECT 108.6000 108.8000 109.0000 109.2000 ;
	    RECT 107.8000 108.2000 108.1000 108.8000 ;
	    RECT 108.6000 108.2000 108.9000 108.8000 ;
	    RECT 107.8000 107.8000 108.2000 108.2000 ;
	    RECT 108.6000 107.8000 109.0000 108.2000 ;
	    RECT 109.4000 105.8000 109.8000 106.2000 ;
	    RECT 109.4000 105.2000 109.7000 105.8000 ;
	    RECT 109.4000 104.8000 109.8000 105.2000 ;
	    RECT 111.0000 103.1000 111.3000 111.8000 ;
	    RECT 112.6000 107.2000 112.9000 113.8000 ;
	    RECT 113.4000 112.1000 113.8000 117.9000 ;
	    RECT 115.0000 114.8000 115.4000 115.2000 ;
	    RECT 116.6000 115.1000 117.0000 115.2000 ;
	    RECT 117.4000 115.1000 117.8000 115.2000 ;
	    RECT 116.6000 114.8000 117.8000 115.1000 ;
	    RECT 115.0000 114.2000 115.3000 114.8000 ;
	    RECT 115.0000 113.8000 115.4000 114.2000 ;
	    RECT 118.2000 112.1000 118.6000 117.9000 ;
	    RECT 123.8000 113.8000 124.2000 114.2000 ;
	    RECT 120.6000 111.8000 121.0000 112.2000 ;
	    RECT 114.2000 110.8000 114.6000 111.2000 ;
	    RECT 113.4000 109.8000 113.8000 110.2000 ;
	    RECT 112.6000 106.8000 113.0000 107.2000 ;
	    RECT 113.4000 106.2000 113.7000 109.8000 ;
	    RECT 113.4000 105.8000 113.8000 106.2000 ;
	    RECT 111.0000 102.8000 112.1000 103.1000 ;
	    RECT 111.0000 101.8000 111.4000 102.2000 ;
	    RECT 108.6000 94.7000 109.0000 95.1000 ;
	    RECT 108.6000 89.2000 108.9000 94.7000 ;
	    RECT 109.4000 92.1000 109.8000 97.9000 ;
	    RECT 111.0000 97.2000 111.3000 101.8000 ;
	    RECT 111.0000 96.8000 111.4000 97.2000 ;
	    RECT 111.8000 96.2000 112.1000 102.8000 ;
	    RECT 111.0000 93.1000 111.4000 95.9000 ;
	    RECT 111.8000 95.8000 112.2000 96.2000 ;
	    RECT 113.4000 95.2000 113.7000 105.8000 ;
	    RECT 114.2000 105.2000 114.5000 110.8000 ;
	    RECT 120.6000 108.2000 120.9000 111.8000 ;
	    RECT 123.8000 109.2000 124.1000 113.8000 ;
	    RECT 128.6000 112.1000 129.0000 117.9000 ;
	    RECT 129.4000 114.8000 129.8000 115.2000 ;
	    RECT 129.4000 114.2000 129.7000 114.8000 ;
	    RECT 132.6000 114.7000 133.0000 115.1000 ;
	    RECT 129.4000 113.8000 129.8000 114.2000 ;
	    RECT 129.4000 112.8000 129.8000 113.2000 ;
	    RECT 129.4000 109.2000 129.7000 112.8000 ;
	    RECT 132.6000 109.2000 132.9000 114.7000 ;
	    RECT 133.4000 112.1000 133.8000 117.9000 ;
	    RECT 135.0000 113.1000 135.4000 115.9000 ;
	    RECT 135.8000 114.8000 136.2000 115.2000 ;
	    RECT 140.6000 115.1000 141.0000 115.2000 ;
	    RECT 141.4000 115.1000 141.8000 115.2000 ;
	    RECT 140.6000 114.8000 141.8000 115.1000 ;
	    RECT 143.0000 115.1000 143.4000 115.2000 ;
	    RECT 143.8000 115.1000 144.2000 115.2000 ;
	    RECT 143.0000 114.8000 144.2000 115.1000 ;
	    RECT 144.6000 115.1000 145.0000 115.2000 ;
	    RECT 145.4000 115.1000 145.8000 115.2000 ;
	    RECT 144.6000 114.8000 145.8000 115.1000 ;
	    RECT 135.8000 109.2000 136.1000 114.8000 ;
	    RECT 139.8000 113.8000 140.2000 114.2000 ;
	    RECT 123.8000 108.8000 124.2000 109.2000 ;
	    RECT 129.4000 108.8000 129.8000 109.2000 ;
	    RECT 132.6000 108.8000 133.0000 109.2000 ;
	    RECT 134.2000 108.8000 134.6000 109.2000 ;
	    RECT 135.8000 108.8000 136.2000 109.2000 ;
	    RECT 134.2000 108.2000 134.5000 108.8000 ;
	    RECT 116.6000 107.8000 117.0000 108.2000 ;
	    RECT 120.6000 107.8000 121.0000 108.2000 ;
	    RECT 124.6000 108.1000 125.0000 108.2000 ;
	    RECT 125.4000 108.1000 125.8000 108.2000 ;
	    RECT 124.6000 107.8000 125.8000 108.1000 ;
	    RECT 134.2000 107.8000 134.6000 108.2000 ;
	    RECT 138.2000 107.8000 138.6000 108.2000 ;
	    RECT 116.6000 107.2000 116.9000 107.8000 ;
	    RECT 138.2000 107.2000 138.5000 107.8000 ;
	    RECT 116.6000 106.8000 117.0000 107.2000 ;
	    RECT 121.4000 106.8000 121.8000 107.2000 ;
	    RECT 122.2000 106.8000 122.6000 107.2000 ;
	    RECT 127.8000 107.1000 128.2000 107.2000 ;
	    RECT 128.6000 107.1000 129.0000 107.2000 ;
	    RECT 127.8000 106.8000 129.0000 107.1000 ;
	    RECT 131.0000 106.8000 131.4000 107.2000 ;
	    RECT 131.8000 106.8000 132.2000 107.2000 ;
	    RECT 138.2000 106.8000 138.6000 107.2000 ;
	    RECT 115.8000 106.1000 116.2000 106.2000 ;
	    RECT 116.6000 106.1000 117.0000 106.2000 ;
	    RECT 115.8000 105.8000 117.0000 106.1000 ;
	    RECT 117.4000 105.8000 117.8000 106.2000 ;
	    RECT 120.6000 105.8000 121.0000 106.2000 ;
	    RECT 117.4000 105.2000 117.7000 105.8000 ;
	    RECT 114.2000 104.8000 114.6000 105.2000 ;
	    RECT 117.4000 104.8000 117.8000 105.2000 ;
	    RECT 120.6000 104.2000 120.9000 105.8000 ;
	    RECT 121.4000 105.2000 121.7000 106.8000 ;
	    RECT 122.2000 106.2000 122.5000 106.8000 ;
	    RECT 131.0000 106.2000 131.3000 106.8000 ;
	    RECT 122.2000 105.8000 122.6000 106.2000 ;
	    RECT 127.0000 105.8000 127.4000 106.2000 ;
	    RECT 128.6000 106.1000 129.0000 106.2000 ;
	    RECT 129.4000 106.1000 129.8000 106.2000 ;
	    RECT 128.6000 105.8000 129.8000 106.1000 ;
	    RECT 131.0000 105.8000 131.4000 106.2000 ;
	    RECT 127.0000 105.2000 127.3000 105.8000 ;
	    RECT 121.4000 104.8000 121.8000 105.2000 ;
	    RECT 127.0000 104.8000 127.4000 105.2000 ;
	    RECT 130.2000 104.8000 130.6000 105.2000 ;
	    RECT 130.2000 104.2000 130.5000 104.8000 ;
	    RECT 120.6000 103.8000 121.0000 104.2000 ;
	    RECT 128.6000 103.8000 129.0000 104.2000 ;
	    RECT 130.2000 103.8000 130.6000 104.2000 ;
	    RECT 128.6000 103.2000 128.9000 103.8000 ;
	    RECT 128.6000 102.8000 129.0000 103.2000 ;
	    RECT 119.0000 101.8000 119.4000 102.2000 ;
	    RECT 119.0000 97.2000 119.3000 101.8000 ;
	    RECT 125.4000 97.8000 125.8000 98.2000 ;
	    RECT 125.4000 97.2000 125.7000 97.8000 ;
	    RECT 115.8000 96.8000 116.2000 97.2000 ;
	    RECT 119.0000 96.8000 119.4000 97.2000 ;
	    RECT 123.8000 96.8000 124.2000 97.2000 ;
	    RECT 125.4000 96.8000 125.8000 97.2000 ;
	    RECT 115.0000 95.8000 115.4000 96.2000 ;
	    RECT 115.0000 95.2000 115.3000 95.8000 ;
	    RECT 113.4000 94.8000 113.8000 95.2000 ;
	    RECT 115.0000 94.8000 115.4000 95.2000 ;
	    RECT 112.6000 94.1000 113.0000 94.2000 ;
	    RECT 113.4000 94.1000 113.8000 94.2000 ;
	    RECT 112.6000 93.8000 113.8000 94.1000 ;
	    RECT 114.2000 93.8000 114.6000 94.2000 ;
	    RECT 114.2000 90.2000 114.5000 93.8000 ;
	    RECT 115.0000 91.2000 115.3000 94.8000 ;
	    RECT 115.0000 90.8000 115.4000 91.2000 ;
	    RECT 114.2000 89.8000 114.6000 90.2000 ;
	    RECT 108.6000 88.8000 109.0000 89.2000 ;
	    RECT 114.2000 89.1000 114.6000 89.2000 ;
	    RECT 115.0000 89.1000 115.4000 89.2000 ;
	    RECT 114.2000 88.8000 115.4000 89.1000 ;
	    RECT 107.0000 86.8000 107.4000 87.2000 ;
	    RECT 109.4000 87.1000 109.8000 87.2000 ;
	    RECT 110.2000 87.1000 110.6000 87.2000 ;
	    RECT 109.4000 86.8000 110.6000 87.1000 ;
	    RECT 107.0000 84.2000 107.3000 86.8000 ;
	    RECT 115.8000 86.2000 116.1000 96.8000 ;
	    RECT 123.8000 96.2000 124.1000 96.8000 ;
	    RECT 116.6000 95.8000 117.0000 96.2000 ;
	    RECT 117.4000 95.8000 117.8000 96.2000 ;
	    RECT 119.0000 95.8000 119.4000 96.2000 ;
	    RECT 123.8000 95.8000 124.2000 96.2000 ;
	    RECT 127.0000 95.8000 127.4000 96.2000 ;
	    RECT 116.6000 95.2000 116.9000 95.8000 ;
	    RECT 117.4000 95.2000 117.7000 95.8000 ;
	    RECT 119.0000 95.2000 119.3000 95.8000 ;
	    RECT 116.6000 94.8000 117.0000 95.2000 ;
	    RECT 117.4000 94.8000 117.8000 95.2000 ;
	    RECT 119.0000 94.8000 119.4000 95.2000 ;
	    RECT 121.4000 95.1000 121.8000 95.2000 ;
	    RECT 122.2000 95.1000 122.6000 95.2000 ;
	    RECT 121.4000 94.8000 122.6000 95.1000 ;
	    RECT 125.4000 95.1000 125.8000 95.2000 ;
	    RECT 126.2000 95.1000 126.6000 95.2000 ;
	    RECT 125.4000 94.8000 126.6000 95.1000 ;
	    RECT 117.4000 93.8000 117.8000 94.2000 ;
	    RECT 117.4000 92.2000 117.7000 93.8000 ;
	    RECT 117.4000 91.8000 117.8000 92.2000 ;
	    RECT 116.6000 90.8000 117.0000 91.2000 ;
	    RECT 116.6000 87.2000 116.9000 90.8000 ;
	    RECT 119.0000 87.2000 119.3000 94.8000 ;
	    RECT 123.8000 94.1000 124.2000 94.2000 ;
	    RECT 124.6000 94.1000 125.0000 94.2000 ;
	    RECT 123.8000 93.8000 125.0000 94.1000 ;
	    RECT 125.4000 93.2000 125.7000 94.8000 ;
	    RECT 127.0000 94.2000 127.3000 95.8000 ;
	    RECT 127.0000 93.8000 127.4000 94.2000 ;
	    RECT 125.4000 92.8000 125.8000 93.2000 ;
	    RECT 127.8000 93.1000 128.2000 95.9000 ;
	    RECT 123.8000 92.1000 124.2000 92.2000 ;
	    RECT 124.6000 92.1000 125.0000 92.2000 ;
	    RECT 129.4000 92.1000 129.8000 97.9000 ;
	    RECT 130.2000 94.7000 130.6000 95.1000 ;
	    RECT 130.2000 92.2000 130.5000 94.7000 ;
	    RECT 123.8000 91.8000 125.0000 92.1000 ;
	    RECT 130.2000 91.8000 130.6000 92.2000 ;
	    RECT 121.4000 89.8000 121.8000 90.2000 ;
	    RECT 121.4000 89.2000 121.7000 89.8000 ;
	    RECT 121.4000 88.8000 121.8000 89.2000 ;
	    RECT 116.6000 86.8000 117.0000 87.2000 ;
	    RECT 119.0000 86.8000 119.4000 87.2000 ;
	    RECT 119.8000 87.1000 120.2000 87.2000 ;
	    RECT 120.6000 87.1000 121.0000 87.2000 ;
	    RECT 119.8000 86.8000 121.0000 87.1000 ;
	    RECT 107.8000 86.1000 108.2000 86.2000 ;
	    RECT 108.6000 86.1000 109.0000 86.2000 ;
	    RECT 107.8000 85.8000 109.0000 86.1000 ;
	    RECT 110.2000 86.1000 110.6000 86.2000 ;
	    RECT 111.0000 86.1000 111.4000 86.2000 ;
	    RECT 110.2000 85.8000 111.4000 86.1000 ;
	    RECT 114.2000 85.8000 114.6000 86.2000 ;
	    RECT 115.8000 85.8000 116.2000 86.2000 ;
	    RECT 108.4000 85.1000 108.8000 85.2000 ;
	    RECT 109.4000 85.1000 109.8000 85.2000 ;
	    RECT 110.2000 85.1000 110.6000 85.2000 ;
	    RECT 108.4000 84.8000 108.9000 85.1000 ;
	    RECT 109.4000 84.8000 110.6000 85.1000 ;
	    RECT 108.6000 84.2000 108.9000 84.8000 ;
	    RECT 114.2000 84.2000 114.5000 85.8000 ;
	    RECT 116.6000 85.2000 116.9000 86.8000 ;
	    RECT 119.0000 86.2000 119.3000 86.8000 ;
	    RECT 119.0000 85.8000 119.4000 86.2000 ;
	    RECT 116.6000 84.8000 117.0000 85.2000 ;
	    RECT 119.8000 84.8000 120.2000 85.2000 ;
	    RECT 107.0000 83.8000 107.4000 84.2000 ;
	    RECT 108.6000 83.8000 109.0000 84.2000 ;
	    RECT 114.2000 83.8000 114.6000 84.2000 ;
	    RECT 106.2000 81.8000 106.6000 82.2000 ;
	    RECT 103.8000 77.8000 104.2000 78.2000 ;
	    RECT 103.8000 75.8000 104.2000 76.2000 ;
	    RECT 103.8000 75.2000 104.1000 75.8000 ;
	    RECT 103.8000 74.8000 104.2000 75.2000 ;
	    RECT 103.8000 74.2000 104.1000 74.8000 ;
	    RECT 106.2000 74.2000 106.5000 81.8000 ;
	    RECT 109.4000 79.8000 109.8000 80.2000 ;
	    RECT 108.6000 77.8000 109.0000 78.2000 ;
	    RECT 108.6000 77.2000 108.9000 77.8000 ;
	    RECT 107.0000 77.1000 107.4000 77.2000 ;
	    RECT 107.8000 77.1000 108.2000 77.2000 ;
	    RECT 107.0000 76.8000 108.2000 77.1000 ;
	    RECT 108.6000 76.8000 109.0000 77.2000 ;
	    RECT 109.4000 76.2000 109.7000 79.8000 ;
	    RECT 110.2000 78.8000 110.6000 79.2000 ;
	    RECT 109.4000 75.8000 109.8000 76.2000 ;
	    RECT 108.6000 74.8000 109.0000 75.2000 ;
	    RECT 103.8000 73.8000 104.2000 74.2000 ;
	    RECT 104.6000 73.8000 105.0000 74.2000 ;
	    RECT 106.2000 73.8000 106.6000 74.2000 ;
	    RECT 99.8000 68.8000 100.2000 69.2000 ;
	    RECT 100.6000 68.8000 101.0000 69.2000 ;
	    RECT 100.6000 68.2000 100.9000 68.8000 ;
	    RECT 100.6000 67.8000 101.0000 68.2000 ;
	    RECT 103.0000 66.1000 103.4000 66.2000 ;
	    RECT 103.8000 66.1000 104.1000 73.8000 ;
	    RECT 104.6000 67.2000 104.9000 73.8000 ;
	    RECT 105.4000 72.8000 105.8000 73.2000 ;
	    RECT 105.4000 71.2000 105.7000 72.8000 ;
	    RECT 105.4000 70.8000 105.8000 71.2000 ;
	    RECT 105.4000 68.2000 105.7000 70.8000 ;
	    RECT 105.4000 67.8000 105.8000 68.2000 ;
	    RECT 106.2000 67.2000 106.5000 73.8000 ;
	    RECT 108.6000 73.2000 108.9000 74.8000 ;
	    RECT 108.6000 72.8000 109.0000 73.2000 ;
	    RECT 104.6000 66.8000 105.0000 67.2000 ;
	    RECT 106.2000 66.8000 106.6000 67.2000 ;
	    RECT 109.4000 67.1000 109.7000 75.8000 ;
	    RECT 110.2000 74.2000 110.5000 78.8000 ;
	    RECT 114.2000 77.8000 114.6000 78.2000 ;
	    RECT 114.2000 77.2000 114.5000 77.8000 ;
	    RECT 114.2000 76.8000 114.6000 77.2000 ;
	    RECT 116.6000 76.2000 116.9000 84.8000 ;
	    RECT 119.8000 84.2000 120.1000 84.8000 ;
	    RECT 118.2000 83.8000 118.6000 84.2000 ;
	    RECT 119.8000 83.8000 120.2000 84.2000 ;
	    RECT 120.6000 83.8000 121.0000 84.2000 ;
	    RECT 118.2000 83.2000 118.5000 83.8000 ;
	    RECT 118.2000 82.8000 118.6000 83.2000 ;
	    RECT 119.0000 81.8000 119.4000 82.2000 ;
	    RECT 111.8000 75.8000 112.2000 76.2000 ;
	    RECT 112.6000 75.8000 113.0000 76.2000 ;
	    RECT 115.8000 76.1000 116.2000 76.2000 ;
	    RECT 115.0000 75.8000 116.2000 76.1000 ;
	    RECT 116.6000 75.8000 117.0000 76.2000 ;
	    RECT 111.8000 75.2000 112.1000 75.8000 ;
	    RECT 111.8000 74.8000 112.2000 75.2000 ;
	    RECT 110.2000 73.8000 110.6000 74.2000 ;
	    RECT 112.6000 70.2000 112.9000 75.8000 ;
	    RECT 113.4000 75.1000 113.8000 75.2000 ;
	    RECT 114.2000 75.1000 114.6000 75.2000 ;
	    RECT 113.4000 74.8000 114.6000 75.1000 ;
	    RECT 113.4000 73.8000 113.8000 74.2000 ;
	    RECT 113.4000 72.2000 113.7000 73.8000 ;
	    RECT 114.2000 72.8000 114.6000 73.2000 ;
	    RECT 113.4000 71.8000 113.8000 72.2000 ;
	    RECT 112.6000 69.8000 113.0000 70.2000 ;
	    RECT 108.6000 66.8000 109.7000 67.1000 ;
	    RECT 110.2000 66.8000 110.6000 67.2000 ;
	    RECT 111.8000 67.1000 112.2000 67.2000 ;
	    RECT 112.6000 67.1000 113.0000 67.2000 ;
	    RECT 111.8000 66.8000 113.0000 67.1000 ;
	    RECT 108.6000 66.2000 108.9000 66.8000 ;
	    RECT 103.0000 65.8000 104.1000 66.1000 ;
	    RECT 104.6000 66.1000 105.0000 66.2000 ;
	    RECT 105.4000 66.1000 105.8000 66.2000 ;
	    RECT 104.6000 65.8000 105.8000 66.1000 ;
	    RECT 108.6000 65.8000 109.0000 66.2000 ;
	    RECT 109.4000 65.8000 109.8000 66.2000 ;
	    RECT 103.8000 65.2000 104.1000 65.8000 ;
	    RECT 103.8000 64.8000 104.2000 65.2000 ;
	    RECT 107.8000 64.8000 108.2000 65.2000 ;
	    RECT 94.2000 62.8000 94.6000 63.2000 ;
	    RECT 96.6000 62.8000 97.0000 63.2000 ;
	    RECT 91.8000 57.8000 92.2000 58.2000 ;
	    RECT 80.6000 54.8000 81.0000 55.2000 ;
	    RECT 81.4000 55.1000 81.8000 55.2000 ;
	    RECT 82.2000 55.1000 82.6000 55.2000 ;
	    RECT 81.4000 54.8000 82.6000 55.1000 ;
	    RECT 86.2000 54.8000 86.6000 55.2000 ;
	    RECT 90.2000 54.8000 90.6000 55.2000 ;
	    RECT 91.0000 54.8000 91.4000 55.2000 ;
	    RECT 79.8000 51.8000 80.2000 52.2000 ;
	    RECT 80.6000 50.2000 80.9000 54.8000 ;
	    RECT 81.4000 53.8000 81.8000 54.2000 ;
	    RECT 81.4000 52.2000 81.7000 53.8000 ;
	    RECT 82.2000 52.2000 82.5000 54.8000 ;
	    RECT 87.0000 53.8000 87.4000 54.2000 ;
	    RECT 87.0000 53.2000 87.3000 53.8000 ;
	    RECT 90.2000 53.2000 90.5000 54.8000 ;
	    RECT 91.8000 54.2000 92.1000 57.8000 ;
	    RECT 94.2000 57.2000 94.5000 62.8000 ;
	    RECT 103.8000 60.2000 104.1000 64.8000 ;
	    RECT 107.8000 64.2000 108.1000 64.8000 ;
	    RECT 106.2000 63.8000 106.6000 64.2000 ;
	    RECT 107.8000 63.8000 108.2000 64.2000 ;
	    RECT 96.6000 59.8000 97.0000 60.2000 ;
	    RECT 103.8000 59.8000 104.2000 60.2000 ;
	    RECT 96.6000 59.2000 96.9000 59.8000 ;
	    RECT 96.6000 58.8000 97.0000 59.2000 ;
	    RECT 103.0000 58.8000 103.4000 59.2000 ;
	    RECT 94.2000 56.8000 94.6000 57.2000 ;
	    RECT 92.6000 55.8000 93.0000 56.2000 ;
	    RECT 92.6000 55.2000 92.9000 55.8000 ;
	    RECT 94.2000 55.2000 94.5000 56.8000 ;
	    RECT 92.6000 54.8000 93.0000 55.2000 ;
	    RECT 94.2000 54.8000 94.6000 55.2000 ;
	    RECT 91.8000 53.8000 92.2000 54.2000 ;
	    RECT 93.4000 53.8000 93.8000 54.2000 ;
	    RECT 93.4000 53.2000 93.7000 53.8000 ;
	    RECT 87.0000 52.8000 87.4000 53.2000 ;
	    RECT 90.2000 52.8000 90.6000 53.2000 ;
	    RECT 91.0000 52.8000 91.4000 53.2000 ;
	    RECT 93.4000 52.8000 93.8000 53.2000 ;
	    RECT 87.0000 52.2000 87.3000 52.8000 ;
	    RECT 81.4000 51.8000 81.8000 52.2000 ;
	    RECT 82.2000 51.8000 82.6000 52.2000 ;
	    RECT 83.8000 51.8000 84.2000 52.2000 ;
	    RECT 87.0000 51.8000 87.4000 52.2000 ;
	    RECT 89.4000 52.1000 89.8000 52.2000 ;
	    RECT 90.2000 52.1000 90.6000 52.2000 ;
	    RECT 89.4000 51.8000 90.6000 52.1000 ;
	    RECT 83.0000 50.8000 83.4000 51.2000 ;
	    RECT 83.0000 50.2000 83.3000 50.8000 ;
	    RECT 83.8000 50.2000 84.1000 51.8000 ;
	    RECT 80.6000 49.8000 81.0000 50.2000 ;
	    RECT 83.0000 49.8000 83.4000 50.2000 ;
	    RECT 83.8000 49.8000 84.2000 50.2000 ;
	    RECT 83.0000 49.2000 83.3000 49.8000 ;
	    RECT 79.0000 49.1000 79.4000 49.2000 ;
	    RECT 79.8000 49.1000 80.2000 49.2000 ;
	    RECT 79.0000 48.8000 80.2000 49.1000 ;
	    RECT 82.2000 48.8000 82.6000 49.2000 ;
	    RECT 83.0000 48.8000 83.4000 49.2000 ;
	    RECT 83.8000 48.8000 84.2000 49.2000 ;
	    RECT 82.2000 48.2000 82.5000 48.8000 ;
	    RECT 82.2000 47.8000 82.6000 48.2000 ;
	    RECT 81.4000 46.8000 81.8000 47.2000 ;
	    RECT 79.8000 45.1000 80.2000 45.2000 ;
	    RECT 80.6000 45.1000 81.0000 45.2000 ;
	    RECT 79.8000 44.8000 81.0000 45.1000 ;
	    RECT 81.4000 44.2000 81.7000 46.8000 ;
	    RECT 83.8000 46.2000 84.1000 48.8000 ;
	    RECT 91.0000 47.2000 91.3000 52.8000 ;
	    RECT 99.0000 52.1000 99.4000 57.9000 ;
	    RECT 103.0000 55.1000 103.3000 58.8000 ;
	    RECT 103.0000 54.7000 103.4000 55.1000 ;
	    RECT 100.6000 52.8000 101.0000 53.2000 ;
	    RECT 93.4000 48.8000 93.8000 49.2000 ;
	    RECT 86.2000 46.8000 86.6000 47.2000 ;
	    RECT 89.4000 46.8000 89.8000 47.2000 ;
	    RECT 90.2000 46.8000 90.6000 47.2000 ;
	    RECT 91.0000 46.8000 91.4000 47.2000 ;
	    RECT 86.2000 46.2000 86.5000 46.8000 ;
	    RECT 83.8000 45.8000 84.2000 46.2000 ;
	    RECT 86.2000 45.8000 86.6000 46.2000 ;
	    RECT 83.8000 45.1000 84.2000 45.2000 ;
	    RECT 84.6000 45.1000 85.0000 45.2000 ;
	    RECT 83.8000 44.8000 85.0000 45.1000 ;
	    RECT 81.4000 43.8000 81.8000 44.2000 ;
	    RECT 79.8000 37.8000 80.2000 38.2000 ;
	    RECT 79.8000 37.2000 80.1000 37.8000 ;
	    RECT 79.0000 36.8000 79.4000 37.2000 ;
	    RECT 79.8000 36.8000 80.2000 37.2000 ;
	    RECT 83.0000 36.8000 83.4000 37.2000 ;
	    RECT 74.2000 34.8000 74.6000 35.2000 ;
	    RECT 75.8000 34.8000 76.2000 35.2000 ;
	    RECT 76.6000 34.8000 77.0000 35.2000 ;
	    RECT 78.2000 34.8000 78.6000 35.2000 ;
	    RECT 74.2000 34.2000 74.5000 34.8000 ;
	    RECT 75.8000 34.2000 76.1000 34.8000 ;
	    RECT 74.2000 33.8000 74.6000 34.2000 ;
	    RECT 75.8000 33.8000 76.2000 34.2000 ;
	    RECT 72.6000 29.8000 73.0000 30.2000 ;
	    RECT 67.8000 26.8000 68.2000 27.2000 ;
	    RECT 71.8000 26.8000 72.2000 27.2000 ;
	    RECT 59.0000 26.1000 59.4000 26.2000 ;
	    RECT 58.2000 25.8000 59.4000 26.1000 ;
	    RECT 47.8000 23.8000 48.2000 24.2000 ;
	    RECT 47.8000 23.2000 48.1000 23.8000 ;
	    RECT 48.6000 23.2000 48.9000 25.8000 ;
	    RECT 50.2000 25.2000 50.5000 25.8000 ;
	    RECT 50.2000 24.8000 50.6000 25.2000 ;
	    RECT 49.4000 23.8000 49.8000 24.2000 ;
	    RECT 47.8000 22.8000 48.2000 23.2000 ;
	    RECT 48.6000 22.8000 49.0000 23.2000 ;
	    RECT 48.6000 22.2000 48.9000 22.8000 ;
	    RECT 48.6000 21.8000 49.0000 22.2000 ;
	    RECT 49.4000 14.2000 49.7000 23.8000 ;
	    RECT 45.4000 13.8000 45.8000 14.2000 ;
	    RECT 49.4000 13.8000 49.8000 14.2000 ;
	    RECT 45.4000 13.2000 45.7000 13.8000 ;
	    RECT 45.4000 12.8000 45.8000 13.2000 ;
	    RECT 43.8000 11.8000 44.2000 12.2000 ;
	    RECT 40.6000 10.8000 41.0000 11.2000 ;
	    RECT 43.0000 10.8000 43.4000 11.2000 ;
	    RECT 43.0000 9.2000 43.3000 10.8000 ;
	    RECT 43.8000 10.2000 44.1000 11.8000 ;
	    RECT 51.0000 11.2000 51.3000 25.8000 ;
	    RECT 51.8000 25.2000 52.1000 25.8000 ;
	    RECT 59.8000 25.2000 60.1000 26.8000 ;
	    RECT 60.6000 26.2000 60.9000 26.8000 ;
	    RECT 72.6000 26.2000 72.9000 29.8000 ;
	    RECT 76.6000 28.2000 76.9000 34.8000 ;
	    RECT 79.0000 28.2000 79.3000 36.8000 ;
	    RECT 79.8000 35.2000 80.1000 36.8000 ;
	    RECT 79.8000 34.8000 80.2000 35.2000 ;
	    RECT 83.0000 33.2000 83.3000 36.8000 ;
	    RECT 84.6000 35.8000 85.0000 36.2000 ;
	    RECT 85.4000 35.8000 85.8000 36.2000 ;
	    RECT 84.6000 35.2000 84.9000 35.8000 ;
	    RECT 84.6000 34.8000 85.0000 35.2000 ;
	    RECT 85.4000 34.1000 85.7000 35.8000 ;
	    RECT 84.6000 33.8000 85.7000 34.1000 ;
	    RECT 83.0000 32.8000 83.4000 33.2000 ;
	    RECT 81.4000 31.8000 81.8000 32.2000 ;
	    RECT 81.4000 29.2000 81.7000 31.8000 ;
	    RECT 81.4000 28.8000 81.8000 29.2000 ;
	    RECT 75.8000 27.8000 76.2000 28.2000 ;
	    RECT 76.6000 27.8000 77.0000 28.2000 ;
	    RECT 79.0000 27.8000 79.4000 28.2000 ;
	    RECT 79.8000 27.8000 80.2000 28.2000 ;
	    RECT 75.8000 26.2000 76.1000 27.8000 ;
	    RECT 76.6000 27.2000 76.9000 27.8000 ;
	    RECT 76.6000 26.8000 77.0000 27.2000 ;
	    RECT 60.6000 25.8000 61.0000 26.2000 ;
	    RECT 61.4000 25.8000 61.8000 26.2000 ;
	    RECT 63.8000 26.1000 64.2000 26.2000 ;
	    RECT 64.6000 26.1000 65.0000 26.2000 ;
	    RECT 63.8000 25.8000 65.0000 26.1000 ;
	    RECT 68.6000 25.8000 69.0000 26.2000 ;
	    RECT 72.6000 25.8000 73.0000 26.2000 ;
	    RECT 75.8000 25.8000 76.2000 26.2000 ;
	    RECT 76.6000 25.8000 77.0000 26.2000 ;
	    RECT 51.8000 24.8000 52.2000 25.2000 ;
	    RECT 56.6000 25.1000 57.0000 25.2000 ;
	    RECT 56.6000 24.8000 57.7000 25.1000 ;
	    RECT 57.4000 24.2000 57.7000 24.8000 ;
	    RECT 58.2000 24.8000 58.6000 25.2000 ;
	    RECT 59.8000 24.8000 60.2000 25.2000 ;
	    RECT 55.0000 24.1000 55.4000 24.2000 ;
	    RECT 55.8000 24.1000 56.2000 24.2000 ;
	    RECT 55.0000 23.8000 56.2000 24.1000 ;
	    RECT 57.4000 23.8000 57.8000 24.2000 ;
	    RECT 55.0000 22.8000 55.4000 23.2000 ;
	    RECT 55.0000 19.2000 55.3000 22.8000 ;
	    RECT 51.8000 18.8000 52.2000 19.2000 ;
	    RECT 55.0000 18.8000 55.4000 19.2000 ;
	    RECT 51.8000 15.2000 52.1000 18.8000 ;
	    RECT 52.6000 17.8000 53.0000 18.2000 ;
	    RECT 55.0000 17.8000 55.4000 18.2000 ;
	    RECT 51.8000 14.8000 52.2000 15.2000 ;
	    RECT 52.6000 14.2000 52.9000 17.8000 ;
	    RECT 53.4000 16.1000 53.8000 16.2000 ;
	    RECT 54.2000 16.1000 54.6000 16.2000 ;
	    RECT 53.4000 15.8000 54.6000 16.1000 ;
	    RECT 52.6000 13.8000 53.0000 14.2000 ;
	    RECT 55.0000 14.1000 55.3000 17.8000 ;
	    RECT 57.4000 16.8000 57.8000 17.2000 ;
	    RECT 57.4000 16.2000 57.7000 16.8000 ;
	    RECT 57.4000 15.8000 57.8000 16.2000 ;
	    RECT 55.8000 14.1000 56.2000 14.2000 ;
	    RECT 55.0000 13.8000 56.2000 14.1000 ;
	    RECT 52.6000 13.2000 52.9000 13.8000 ;
	    RECT 51.8000 12.8000 52.2000 13.2000 ;
	    RECT 52.6000 12.8000 53.0000 13.2000 ;
	    RECT 51.8000 12.2000 52.1000 12.8000 ;
	    RECT 51.8000 11.8000 52.2000 12.2000 ;
	    RECT 49.4000 10.8000 49.8000 11.2000 ;
	    RECT 51.0000 10.8000 51.4000 11.2000 ;
	    RECT 43.8000 9.8000 44.2000 10.2000 ;
	    RECT 43.0000 8.8000 43.4000 9.2000 ;
	    RECT 47.0000 8.8000 47.4000 9.2000 ;
	    RECT 47.0000 8.2000 47.3000 8.8000 ;
	    RECT 47.0000 7.8000 47.4000 8.2000 ;
	    RECT 43.8000 6.8000 44.2000 7.2000 ;
	    RECT 38.2000 5.8000 39.3000 6.1000 ;
	    RECT 42.2000 6.1000 42.6000 6.2000 ;
	    RECT 43.0000 6.1000 43.4000 6.2000 ;
	    RECT 42.2000 5.8000 43.4000 6.1000 ;
	    RECT 32.6000 5.2000 32.9000 5.8000 ;
	    RECT 43.8000 5.2000 44.1000 6.8000 ;
	    RECT 47.0000 6.2000 47.3000 7.8000 ;
	    RECT 49.4000 7.2000 49.7000 10.8000 ;
	    RECT 48.6000 7.1000 49.0000 7.2000 ;
	    RECT 49.4000 7.1000 49.8000 7.2000 ;
	    RECT 48.6000 6.8000 49.8000 7.1000 ;
	    RECT 52.6000 6.2000 52.9000 12.8000 ;
	    RECT 55.8000 11.8000 56.2000 12.2000 ;
	    RECT 55.8000 9.2000 56.1000 11.8000 ;
	    RECT 53.4000 8.8000 53.8000 9.2000 ;
	    RECT 55.8000 8.8000 56.2000 9.2000 ;
	    RECT 53.4000 8.2000 53.7000 8.8000 ;
	    RECT 53.4000 7.8000 53.8000 8.2000 ;
	    RECT 55.0000 7.8000 55.4000 8.2000 ;
	    RECT 53.4000 6.8000 53.8000 7.2000 ;
	    RECT 53.4000 6.2000 53.7000 6.8000 ;
	    RECT 55.0000 6.2000 55.3000 7.8000 ;
	    RECT 58.2000 7.2000 58.5000 24.8000 ;
	    RECT 59.0000 18.8000 59.4000 19.2000 ;
	    RECT 59.0000 17.2000 59.3000 18.8000 ;
	    RECT 60.6000 17.2000 60.9000 25.8000 ;
	    RECT 61.4000 25.2000 61.7000 25.8000 ;
	    RECT 68.6000 25.2000 68.9000 25.8000 ;
	    RECT 61.4000 24.8000 61.8000 25.2000 ;
	    RECT 65.4000 24.8000 65.8000 25.2000 ;
	    RECT 68.6000 24.8000 69.0000 25.2000 ;
	    RECT 75.8000 25.1000 76.2000 25.2000 ;
	    RECT 76.6000 25.1000 76.9000 25.8000 ;
	    RECT 75.8000 24.8000 76.9000 25.1000 ;
	    RECT 79.0000 25.2000 79.3000 27.8000 ;
	    RECT 79.8000 27.2000 80.1000 27.8000 ;
	    RECT 79.8000 26.8000 80.2000 27.2000 ;
	    RECT 79.0000 24.8000 79.4000 25.2000 ;
	    RECT 65.4000 24.2000 65.7000 24.8000 ;
	    RECT 61.4000 23.8000 61.8000 24.2000 ;
	    RECT 63.0000 24.1000 63.4000 24.2000 ;
	    RECT 63.8000 24.1000 64.2000 24.2000 ;
	    RECT 63.0000 23.8000 64.2000 24.1000 ;
	    RECT 65.4000 23.8000 65.8000 24.2000 ;
	    RECT 61.4000 19.2000 61.7000 23.8000 ;
	    RECT 64.6000 21.8000 65.0000 22.2000 ;
	    RECT 71.0000 21.8000 71.4000 22.2000 ;
	    RECT 64.6000 21.2000 64.9000 21.8000 ;
	    RECT 64.6000 20.8000 65.0000 21.2000 ;
	    RECT 65.4000 19.8000 65.8000 20.2000 ;
	    RECT 61.4000 18.8000 61.8000 19.2000 ;
	    RECT 63.8000 19.1000 64.2000 19.2000 ;
	    RECT 64.6000 19.1000 65.0000 19.2000 ;
	    RECT 63.8000 18.8000 65.0000 19.1000 ;
	    RECT 59.0000 16.8000 59.4000 17.2000 ;
	    RECT 60.6000 16.8000 61.0000 17.2000 ;
	    RECT 63.0000 16.8000 63.4000 17.2000 ;
	    RECT 59.0000 14.2000 59.3000 16.8000 ;
	    RECT 59.0000 13.8000 59.4000 14.2000 ;
	    RECT 63.0000 13.2000 63.3000 16.8000 ;
	    RECT 65.4000 16.2000 65.7000 19.8000 ;
	    RECT 69.4000 18.8000 69.8000 19.2000 ;
	    RECT 69.4000 18.2000 69.7000 18.8000 ;
	    RECT 69.4000 17.8000 69.8000 18.2000 ;
	    RECT 65.4000 15.8000 65.8000 16.2000 ;
	    RECT 66.2000 15.8000 66.6000 16.2000 ;
	    RECT 66.2000 15.2000 66.5000 15.8000 ;
	    RECT 63.8000 14.8000 64.2000 15.2000 ;
	    RECT 65.4000 15.1000 65.8000 15.2000 ;
	    RECT 64.6000 14.8000 65.8000 15.1000 ;
	    RECT 66.2000 14.8000 66.6000 15.2000 ;
	    RECT 68.6000 14.8000 69.0000 15.2000 ;
	    RECT 63.8000 14.2000 64.1000 14.8000 ;
	    RECT 63.8000 13.8000 64.2000 14.2000 ;
	    RECT 59.8000 13.1000 60.2000 13.2000 ;
	    RECT 60.6000 13.1000 61.0000 13.2000 ;
	    RECT 59.8000 12.8000 61.0000 13.1000 ;
	    RECT 63.0000 12.8000 63.4000 13.2000 ;
	    RECT 58.2000 7.1000 58.6000 7.2000 ;
	    RECT 59.0000 7.1000 59.4000 7.2000 ;
	    RECT 58.2000 6.8000 59.4000 7.1000 ;
	    RECT 62.2000 6.8000 62.6000 7.2000 ;
	    RECT 63.0000 7.1000 63.3000 12.8000 ;
	    RECT 63.8000 7.1000 64.2000 7.2000 ;
	    RECT 63.0000 6.8000 64.2000 7.1000 ;
	    RECT 62.2000 6.2000 62.5000 6.8000 ;
	    RECT 64.6000 6.2000 64.9000 14.8000 ;
	    RECT 68.6000 14.2000 68.9000 14.8000 ;
	    RECT 71.0000 14.2000 71.3000 21.8000 ;
	    RECT 71.8000 15.1000 72.2000 15.2000 ;
	    RECT 72.6000 15.1000 73.0000 15.2000 ;
	    RECT 71.8000 14.8000 73.0000 15.1000 ;
	    RECT 76.6000 15.1000 76.9000 24.8000 ;
	    RECT 77.4000 21.8000 77.8000 22.2000 ;
	    RECT 77.4000 20.2000 77.7000 21.8000 ;
	    RECT 77.4000 19.8000 77.8000 20.2000 ;
	    RECT 77.4000 15.1000 77.8000 15.2000 ;
	    RECT 76.6000 14.8000 77.8000 15.1000 ;
	    RECT 68.6000 13.8000 69.0000 14.2000 ;
	    RECT 71.0000 13.8000 71.4000 14.2000 ;
	    RECT 73.4000 14.1000 73.8000 14.2000 ;
	    RECT 74.2000 14.1000 74.6000 14.2000 ;
	    RECT 73.4000 13.8000 74.6000 14.1000 ;
	    RECT 70.2000 13.1000 70.6000 13.2000 ;
	    RECT 71.0000 13.1000 71.4000 13.2000 ;
	    RECT 70.2000 12.8000 71.4000 13.1000 ;
	    RECT 75.0000 12.8000 75.4000 13.2000 ;
	    RECT 78.2000 13.1000 78.6000 13.2000 ;
	    RECT 79.0000 13.1000 79.4000 13.2000 ;
	    RECT 78.2000 12.8000 79.4000 13.1000 ;
	    RECT 75.0000 12.2000 75.3000 12.8000 ;
	    RECT 74.2000 11.8000 74.6000 12.2000 ;
	    RECT 75.0000 11.8000 75.4000 12.2000 ;
	    RECT 70.2000 9.1000 70.6000 9.2000 ;
	    RECT 71.0000 9.1000 71.4000 9.2000 ;
	    RECT 70.2000 8.8000 71.4000 9.1000 ;
	    RECT 69.4000 6.8000 69.8000 7.2000 ;
	    RECT 69.4000 6.2000 69.7000 6.8000 ;
	    RECT 46.2000 5.8000 46.6000 6.2000 ;
	    RECT 47.0000 5.8000 47.4000 6.2000 ;
	    RECT 52.6000 5.8000 53.0000 6.2000 ;
	    RECT 53.4000 5.8000 53.8000 6.2000 ;
	    RECT 55.0000 5.8000 55.4000 6.2000 ;
	    RECT 58.2000 5.8000 58.6000 6.2000 ;
	    RECT 62.2000 5.8000 62.6000 6.2000 ;
	    RECT 63.8000 5.8000 64.2000 6.2000 ;
	    RECT 64.6000 5.8000 65.0000 6.2000 ;
	    RECT 67.0000 6.1000 67.4000 6.2000 ;
	    RECT 67.8000 6.1000 68.2000 6.2000 ;
	    RECT 67.0000 5.8000 68.2000 6.1000 ;
	    RECT 69.4000 5.8000 69.8000 6.2000 ;
	    RECT 46.2000 5.2000 46.5000 5.8000 ;
	    RECT 58.2000 5.2000 58.5000 5.8000 ;
	    RECT 63.8000 5.2000 64.1000 5.8000 ;
	    RECT 10.2000 4.8000 10.6000 5.2000 ;
	    RECT 15.8000 4.8000 16.2000 5.2000 ;
	    RECT 19.0000 4.8000 19.4000 5.2000 ;
	    RECT 25.4000 4.8000 25.8000 5.2000 ;
	    RECT 30.8000 5.1000 31.2000 5.2000 ;
	    RECT 30.8000 4.8000 31.3000 5.1000 ;
	    RECT 32.6000 4.8000 33.0000 5.2000 ;
	    RECT 43.8000 4.8000 44.2000 5.2000 ;
	    RECT 46.2000 4.8000 46.6000 5.2000 ;
	    RECT 50.8000 5.1000 51.2000 5.2000 ;
	    RECT 51.8000 5.1000 52.2000 5.2000 ;
	    RECT 50.8000 4.8000 52.2000 5.1000 ;
	    RECT 58.2000 4.8000 58.6000 5.2000 ;
	    RECT 62.2000 4.8000 62.6000 5.2000 ;
	    RECT 63.8000 4.8000 64.2000 5.2000 ;
	    RECT 66.2000 5.1000 66.6000 5.2000 ;
	    RECT 67.0000 5.1000 67.4000 5.2000 ;
	    RECT 66.2000 4.8000 67.4000 5.1000 ;
	    RECT 19.0000 4.2000 19.3000 4.8000 ;
	    RECT 31.0000 4.2000 31.3000 4.8000 ;
	    RECT 43.8000 4.2000 44.1000 4.8000 ;
	    RECT 62.2000 4.2000 62.5000 4.8000 ;
	    RECT 19.0000 3.8000 19.4000 4.2000 ;
	    RECT 31.0000 3.8000 31.4000 4.2000 ;
	    RECT 43.8000 3.8000 44.2000 4.2000 ;
	    RECT 62.2000 3.8000 62.6000 4.2000 ;
	    RECT 68.6000 4.1000 69.0000 4.2000 ;
	    RECT 69.4000 4.1000 69.8000 4.2000 ;
	    RECT 68.6000 3.8000 69.8000 4.1000 ;
	    RECT 72.6000 3.1000 73.0000 8.9000 ;
	    RECT 74.2000 4.2000 74.5000 11.8000 ;
	    RECT 79.8000 9.2000 80.1000 26.8000 ;
	    RECT 80.6000 26.1000 81.0000 26.2000 ;
	    RECT 81.4000 26.1000 81.8000 26.2000 ;
	    RECT 80.6000 25.8000 81.8000 26.1000 ;
	    RECT 82.2000 25.8000 82.6000 26.2000 ;
	    RECT 82.2000 25.2000 82.5000 25.8000 ;
	    RECT 84.6000 25.2000 84.9000 33.8000 ;
	    RECT 86.2000 33.2000 86.5000 45.8000 ;
	    RECT 89.4000 45.2000 89.7000 46.8000 ;
	    RECT 90.2000 46.2000 90.5000 46.8000 ;
	    RECT 91.0000 46.2000 91.3000 46.8000 ;
	    RECT 93.4000 46.2000 93.7000 48.8000 ;
	    RECT 96.6000 46.8000 97.0000 47.2000 ;
	    RECT 96.6000 46.2000 96.9000 46.8000 ;
	    RECT 100.6000 46.2000 100.9000 52.8000 ;
	    RECT 103.8000 52.1000 104.2000 57.9000 ;
	    RECT 104.6000 53.8000 105.0000 54.2000 ;
	    RECT 102.2000 50.8000 102.6000 51.2000 ;
	    RECT 102.2000 48.2000 102.5000 50.8000 ;
	    RECT 101.4000 48.1000 101.8000 48.2000 ;
	    RECT 102.2000 48.1000 102.6000 48.2000 ;
	    RECT 101.4000 47.8000 102.6000 48.1000 ;
	    RECT 90.2000 45.8000 90.6000 46.2000 ;
	    RECT 91.0000 45.8000 91.4000 46.2000 ;
	    RECT 93.4000 45.8000 93.8000 46.2000 ;
	    RECT 95.8000 45.8000 96.2000 46.2000 ;
	    RECT 96.6000 45.8000 97.0000 46.2000 ;
	    RECT 99.8000 46.1000 100.2000 46.2000 ;
	    RECT 100.6000 46.1000 101.0000 46.2000 ;
	    RECT 99.8000 45.8000 101.0000 46.1000 ;
	    RECT 95.8000 45.2000 96.1000 45.8000 ;
	    RECT 89.4000 44.8000 89.8000 45.2000 ;
	    RECT 94.2000 44.8000 94.6000 45.2000 ;
	    RECT 95.8000 44.8000 96.2000 45.2000 ;
	    RECT 94.2000 44.2000 94.5000 44.8000 ;
	    RECT 88.6000 43.8000 89.0000 44.2000 ;
	    RECT 92.6000 43.8000 93.0000 44.2000 ;
	    RECT 94.2000 43.8000 94.6000 44.2000 ;
	    RECT 95.8000 43.8000 96.2000 44.2000 ;
	    RECT 88.6000 43.2000 88.9000 43.8000 ;
	    RECT 92.6000 43.2000 92.9000 43.8000 ;
	    RECT 95.8000 43.2000 96.1000 43.8000 ;
	    RECT 88.6000 42.8000 89.0000 43.2000 ;
	    RECT 92.6000 42.8000 93.0000 43.2000 ;
	    RECT 95.8000 42.8000 96.2000 43.2000 ;
	    RECT 94.2000 41.8000 94.6000 42.2000 ;
	    RECT 91.0000 38.8000 91.4000 39.2000 ;
	    RECT 87.8000 34.8000 88.2000 35.2000 ;
	    RECT 89.4000 35.1000 89.8000 35.2000 ;
	    RECT 90.2000 35.1000 90.6000 35.2000 ;
	    RECT 89.4000 34.8000 90.6000 35.1000 ;
	    RECT 87.8000 34.2000 88.1000 34.8000 ;
	    RECT 87.8000 33.8000 88.2000 34.2000 ;
	    RECT 86.2000 32.8000 86.6000 33.2000 ;
	    RECT 87.8000 32.8000 88.2000 33.2000 ;
	    RECT 89.4000 32.8000 89.8000 33.2000 ;
	    RECT 87.8000 29.2000 88.1000 32.8000 ;
	    RECT 87.8000 28.8000 88.2000 29.2000 ;
	    RECT 85.4000 27.1000 85.8000 27.2000 ;
	    RECT 86.2000 27.1000 86.6000 27.2000 ;
	    RECT 85.4000 26.8000 86.6000 27.1000 ;
	    RECT 87.0000 26.8000 87.4000 27.2000 ;
	    RECT 87.0000 26.2000 87.3000 26.8000 ;
	    RECT 87.0000 25.8000 87.4000 26.2000 ;
	    RECT 82.2000 24.8000 82.6000 25.2000 ;
	    RECT 83.8000 25.1000 84.2000 25.2000 ;
	    RECT 84.6000 25.1000 85.0000 25.2000 ;
	    RECT 88.6000 25.1000 89.0000 27.9000 ;
	    RECT 89.4000 27.2000 89.7000 32.8000 ;
	    RECT 89.4000 26.8000 89.8000 27.2000 ;
	    RECT 83.8000 24.8000 85.0000 25.1000 ;
	    RECT 83.0000 21.8000 83.4000 22.2000 ;
	    RECT 83.0000 17.2000 83.3000 21.8000 ;
	    RECT 83.0000 16.8000 83.4000 17.2000 ;
	    RECT 80.6000 15.1000 81.0000 15.2000 ;
	    RECT 81.4000 15.1000 81.8000 15.2000 ;
	    RECT 80.6000 14.8000 81.8000 15.1000 ;
	    RECT 84.6000 14.2000 84.9000 24.8000 ;
	    RECT 87.8000 21.8000 88.2000 22.2000 ;
	    RECT 87.8000 16.2000 88.1000 21.8000 ;
	    RECT 87.8000 15.8000 88.2000 16.2000 ;
	    RECT 85.4000 14.8000 85.8000 15.2000 ;
	    RECT 87.0000 15.1000 87.4000 15.2000 ;
	    RECT 87.8000 15.1000 88.2000 15.2000 ;
	    RECT 87.0000 14.8000 88.2000 15.1000 ;
	    RECT 80.6000 14.1000 81.0000 14.2000 ;
	    RECT 81.4000 14.1000 81.8000 14.2000 ;
	    RECT 80.6000 13.8000 81.8000 14.1000 ;
	    RECT 84.6000 13.8000 85.0000 14.2000 ;
	    RECT 85.4000 13.2000 85.7000 14.8000 ;
	    RECT 89.4000 14.2000 89.7000 26.8000 ;
	    RECT 90.2000 23.1000 90.6000 28.9000 ;
	    RECT 91.0000 15.2000 91.3000 38.8000 ;
	    RECT 94.2000 34.2000 94.5000 41.8000 ;
	    RECT 100.6000 38.2000 100.9000 45.8000 ;
	    RECT 104.6000 44.2000 104.9000 53.8000 ;
	    RECT 105.4000 53.1000 105.8000 55.9000 ;
	    RECT 106.2000 55.2000 106.5000 63.8000 ;
	    RECT 107.8000 62.8000 108.2000 63.2000 ;
	    RECT 106.2000 54.8000 106.6000 55.2000 ;
	    RECT 107.8000 53.2000 108.1000 62.8000 ;
	    RECT 108.6000 56.1000 108.9000 65.8000 ;
	    RECT 109.4000 65.2000 109.7000 65.8000 ;
	    RECT 109.4000 64.8000 109.8000 65.2000 ;
	    RECT 110.2000 63.2000 110.5000 66.8000 ;
	    RECT 111.0000 65.8000 111.4000 66.2000 ;
	    RECT 112.6000 65.8000 113.0000 66.2000 ;
	    RECT 111.0000 64.2000 111.3000 65.8000 ;
	    RECT 112.6000 65.2000 112.9000 65.8000 ;
	    RECT 112.6000 64.8000 113.0000 65.2000 ;
	    RECT 114.2000 64.2000 114.5000 72.8000 ;
	    RECT 115.0000 69.2000 115.3000 75.8000 ;
	    RECT 119.0000 75.2000 119.3000 81.8000 ;
	    RECT 119.8000 77.8000 120.2000 78.2000 ;
	    RECT 115.8000 74.8000 116.2000 75.2000 ;
	    RECT 116.6000 74.8000 117.0000 75.2000 ;
	    RECT 119.0000 74.8000 119.4000 75.2000 ;
	    RECT 115.0000 68.8000 115.4000 69.2000 ;
	    RECT 115.8000 66.2000 116.1000 74.8000 ;
	    RECT 116.6000 73.2000 116.9000 74.8000 ;
	    RECT 119.8000 74.2000 120.1000 77.8000 ;
	    RECT 120.6000 75.2000 120.9000 83.8000 ;
	    RECT 125.4000 83.1000 125.8000 88.9000 ;
	    RECT 129.4000 85.9000 129.8000 86.3000 ;
	    RECT 122.2000 82.1000 122.6000 82.2000 ;
	    RECT 123.0000 82.1000 123.4000 82.2000 ;
	    RECT 122.2000 81.8000 123.4000 82.1000 ;
	    RECT 129.4000 82.1000 129.7000 85.9000 ;
	    RECT 130.2000 83.1000 130.6000 88.9000 ;
	    RECT 131.0000 86.2000 131.3000 105.8000 ;
	    RECT 131.8000 105.2000 132.1000 106.8000 ;
	    RECT 135.8000 105.8000 136.2000 106.2000 ;
	    RECT 137.4000 106.1000 137.8000 106.2000 ;
	    RECT 138.2000 106.1000 138.6000 106.2000 ;
	    RECT 137.4000 105.8000 138.6000 106.1000 ;
	    RECT 135.8000 105.2000 136.1000 105.8000 ;
	    RECT 131.8000 104.8000 132.2000 105.2000 ;
	    RECT 135.8000 104.8000 136.2000 105.2000 ;
	    RECT 139.0000 105.1000 139.4000 107.9000 ;
	    RECT 139.8000 107.2000 140.1000 113.8000 ;
	    RECT 139.8000 106.8000 140.2000 107.2000 ;
	    RECT 139.8000 98.2000 140.1000 106.8000 ;
	    RECT 140.6000 103.1000 141.0000 108.9000 ;
	    RECT 141.4000 106.1000 141.8000 106.2000 ;
	    RECT 142.2000 106.1000 142.6000 106.2000 ;
	    RECT 141.4000 105.8000 142.6000 106.1000 ;
	    RECT 133.4000 97.8000 133.8000 98.2000 ;
	    RECT 133.4000 95.2000 133.7000 97.8000 ;
	    RECT 133.4000 94.8000 133.8000 95.2000 ;
	    RECT 131.0000 85.8000 131.4000 86.2000 ;
	    RECT 131.8000 85.1000 132.2000 87.9000 ;
	    RECT 132.6000 85.1000 133.0000 87.9000 ;
	    RECT 133.4000 87.2000 133.7000 94.8000 ;
	    RECT 134.2000 92.1000 134.6000 97.9000 ;
	    RECT 139.8000 97.8000 140.2000 98.2000 ;
	    RECT 136.6000 97.1000 137.0000 97.2000 ;
	    RECT 137.4000 97.1000 137.8000 97.2000 ;
	    RECT 136.6000 96.8000 137.8000 97.1000 ;
	    RECT 140.6000 96.8000 141.0000 97.2000 ;
	    RECT 136.6000 96.2000 136.9000 96.8000 ;
	    RECT 136.6000 95.8000 137.0000 96.2000 ;
	    RECT 140.6000 95.2000 140.9000 96.8000 ;
	    RECT 144.6000 95.2000 144.9000 114.8000 ;
	    RECT 147.0000 109.1000 147.4000 109.2000 ;
	    RECT 147.8000 109.1000 148.2000 109.2000 ;
	    RECT 145.4000 103.1000 145.8000 108.9000 ;
	    RECT 147.0000 108.8000 148.2000 109.1000 ;
	    RECT 146.2000 103.8000 146.6000 104.2000 ;
	    RECT 139.8000 94.8000 140.2000 95.2000 ;
	    RECT 140.6000 94.8000 141.0000 95.2000 ;
	    RECT 143.0000 94.8000 143.4000 95.2000 ;
	    RECT 144.6000 94.8000 145.0000 95.2000 ;
	    RECT 137.4000 94.1000 137.8000 94.2000 ;
	    RECT 138.2000 94.1000 138.6000 94.2000 ;
	    RECT 137.4000 93.8000 138.6000 94.1000 ;
	    RECT 139.0000 93.8000 139.4000 94.2000 ;
	    RECT 139.0000 93.2000 139.3000 93.8000 ;
	    RECT 137.4000 92.8000 137.8000 93.2000 ;
	    RECT 139.0000 92.8000 139.4000 93.2000 ;
	    RECT 133.4000 86.8000 133.8000 87.2000 ;
	    RECT 132.6000 83.8000 133.0000 84.2000 ;
	    RECT 129.4000 81.8000 130.5000 82.1000 ;
	    RECT 122.2000 76.8000 122.6000 77.2000 ;
	    RECT 120.6000 74.8000 121.0000 75.2000 ;
	    RECT 118.2000 73.8000 118.6000 74.2000 ;
	    RECT 119.0000 73.8000 119.4000 74.2000 ;
	    RECT 119.8000 73.8000 120.2000 74.2000 ;
	    RECT 122.2000 74.1000 122.5000 76.8000 ;
	    RECT 123.0000 75.2000 123.3000 81.8000 ;
	    RECT 129.4000 79.8000 129.8000 80.2000 ;
	    RECT 124.6000 76.8000 125.0000 77.2000 ;
	    RECT 124.6000 76.2000 124.9000 76.8000 ;
	    RECT 124.4000 75.8000 124.9000 76.2000 ;
	    RECT 125.4000 75.8000 125.8000 76.2000 ;
	    RECT 123.0000 74.8000 123.4000 75.2000 ;
	    RECT 123.0000 74.1000 123.4000 74.2000 ;
	    RECT 122.2000 73.8000 123.4000 74.1000 ;
	    RECT 118.2000 73.2000 118.5000 73.8000 ;
	    RECT 116.6000 72.8000 117.0000 73.2000 ;
	    RECT 118.2000 72.8000 118.6000 73.2000 ;
	    RECT 117.4000 71.8000 117.8000 72.2000 ;
	    RECT 117.4000 71.2000 117.7000 71.8000 ;
	    RECT 116.6000 70.8000 117.0000 71.2000 ;
	    RECT 117.4000 70.8000 117.8000 71.2000 ;
	    RECT 116.6000 68.2000 116.9000 70.8000 ;
	    RECT 116.6000 67.8000 117.0000 68.2000 ;
	    RECT 115.0000 65.8000 115.4000 66.2000 ;
	    RECT 115.8000 65.8000 116.2000 66.2000 ;
	    RECT 115.0000 65.2000 115.3000 65.8000 ;
	    RECT 115.8000 65.2000 116.1000 65.8000 ;
	    RECT 115.0000 64.8000 115.4000 65.2000 ;
	    RECT 115.8000 64.8000 116.2000 65.2000 ;
	    RECT 116.6000 64.2000 116.9000 67.8000 ;
	    RECT 117.4000 65.8000 117.8000 66.2000 ;
	    RECT 118.2000 66.1000 118.6000 66.2000 ;
	    RECT 119.0000 66.1000 119.3000 73.8000 ;
	    RECT 123.0000 73.2000 123.3000 73.8000 ;
	    RECT 123.0000 72.8000 123.4000 73.2000 ;
	    RECT 122.2000 71.8000 122.6000 72.2000 ;
	    RECT 122.2000 67.2000 122.5000 71.8000 ;
	    RECT 124.6000 68.8000 125.0000 69.2000 ;
	    RECT 124.6000 68.2000 124.9000 68.8000 ;
	    RECT 124.6000 67.8000 125.0000 68.2000 ;
	    RECT 125.4000 67.2000 125.7000 75.8000 ;
	    RECT 126.2000 75.1000 126.6000 75.2000 ;
	    RECT 127.0000 75.1000 127.4000 75.2000 ;
	    RECT 126.2000 74.8000 127.4000 75.1000 ;
	    RECT 126.2000 73.8000 126.6000 74.2000 ;
	    RECT 126.2000 73.2000 126.5000 73.8000 ;
	    RECT 126.2000 72.8000 126.6000 73.2000 ;
	    RECT 127.0000 68.1000 127.3000 74.8000 ;
	    RECT 129.4000 69.2000 129.7000 79.8000 ;
	    RECT 130.2000 79.2000 130.5000 81.8000 ;
	    RECT 130.2000 78.8000 130.6000 79.2000 ;
	    RECT 130.2000 76.8000 130.6000 77.2000 ;
	    RECT 131.8000 76.8000 132.2000 77.2000 ;
	    RECT 130.2000 75.2000 130.5000 76.8000 ;
	    RECT 131.8000 76.2000 132.1000 76.8000 ;
	    RECT 131.8000 75.8000 132.2000 76.2000 ;
	    RECT 130.2000 74.8000 130.6000 75.2000 ;
	    RECT 132.6000 74.2000 132.9000 83.8000 ;
	    RECT 134.2000 83.1000 134.6000 88.9000 ;
	    RECT 135.0000 85.9000 135.4000 86.3000 ;
	    RECT 135.0000 80.2000 135.3000 85.9000 ;
	    RECT 135.0000 79.8000 135.4000 80.2000 ;
	    RECT 136.6000 75.8000 137.0000 76.2000 ;
	    RECT 136.6000 75.2000 136.9000 75.8000 ;
	    RECT 135.0000 74.8000 135.4000 75.2000 ;
	    RECT 136.6000 74.8000 137.0000 75.2000 ;
	    RECT 132.6000 73.8000 133.0000 74.2000 ;
	    RECT 134.2000 73.8000 134.6000 74.2000 ;
	    RECT 130.2000 72.8000 130.6000 73.2000 ;
	    RECT 129.4000 68.8000 129.8000 69.2000 ;
	    RECT 130.2000 68.2000 130.5000 72.8000 ;
	    RECT 134.2000 72.2000 134.5000 73.8000 ;
	    RECT 135.0000 72.2000 135.3000 74.8000 ;
	    RECT 137.4000 73.2000 137.7000 92.8000 ;
	    RECT 139.0000 83.1000 139.4000 88.9000 ;
	    RECT 138.2000 77.8000 138.6000 78.2000 ;
	    RECT 138.2000 77.2000 138.5000 77.8000 ;
	    RECT 138.2000 76.8000 138.6000 77.2000 ;
	    RECT 139.8000 75.2000 140.1000 94.8000 ;
	    RECT 143.0000 94.2000 143.3000 94.8000 ;
	    RECT 143.0000 93.8000 143.4000 94.2000 ;
	    RECT 144.6000 93.2000 144.9000 94.8000 ;
	    RECT 143.0000 92.8000 143.4000 93.2000 ;
	    RECT 144.6000 92.8000 145.0000 93.2000 ;
	    RECT 143.0000 89.2000 143.3000 92.8000 ;
	    RECT 143.0000 88.8000 143.4000 89.2000 ;
	    RECT 144.6000 85.8000 145.0000 86.2000 ;
	    RECT 145.4000 85.8000 145.8000 86.2000 ;
	    RECT 141.4000 84.1000 141.8000 84.2000 ;
	    RECT 142.2000 84.1000 142.6000 84.2000 ;
	    RECT 141.4000 83.8000 142.6000 84.1000 ;
	    RECT 143.0000 81.8000 143.4000 82.2000 ;
	    RECT 143.0000 77.2000 143.3000 81.8000 ;
	    RECT 144.6000 81.2000 144.9000 85.8000 ;
	    RECT 145.4000 84.2000 145.7000 85.8000 ;
	    RECT 145.4000 83.8000 145.8000 84.2000 ;
	    RECT 144.6000 80.8000 145.0000 81.2000 ;
	    RECT 143.0000 76.8000 143.4000 77.2000 ;
	    RECT 145.4000 76.8000 145.8000 77.2000 ;
	    RECT 138.2000 74.8000 138.6000 75.2000 ;
	    RECT 139.8000 74.8000 140.2000 75.2000 ;
	    RECT 142.2000 75.1000 142.6000 75.2000 ;
	    RECT 143.0000 75.1000 143.4000 75.2000 ;
	    RECT 142.2000 74.8000 143.4000 75.1000 ;
	    RECT 143.8000 74.8000 144.2000 75.2000 ;
	    RECT 137.4000 72.8000 137.8000 73.2000 ;
	    RECT 133.4000 71.8000 133.8000 72.2000 ;
	    RECT 134.2000 71.8000 134.6000 72.2000 ;
	    RECT 135.0000 71.8000 135.4000 72.2000 ;
	    RECT 137.4000 71.8000 137.8000 72.2000 ;
	    RECT 133.4000 71.2000 133.7000 71.8000 ;
	    RECT 133.4000 70.8000 133.8000 71.2000 ;
	    RECT 136.6000 70.8000 137.0000 71.2000 ;
	    RECT 133.4000 70.2000 133.7000 70.8000 ;
	    RECT 133.4000 69.8000 133.8000 70.2000 ;
	    RECT 135.8000 68.8000 136.2000 69.2000 ;
	    RECT 126.2000 67.8000 127.3000 68.1000 ;
	    RECT 127.8000 67.8000 128.2000 68.2000 ;
	    RECT 130.2000 67.8000 130.6000 68.2000 ;
	    RECT 133.4000 67.8000 133.8000 68.2000 ;
	    RECT 126.2000 67.2000 126.5000 67.8000 ;
	    RECT 122.2000 66.8000 122.6000 67.2000 ;
	    RECT 123.0000 66.8000 123.4000 67.2000 ;
	    RECT 124.6000 66.8000 125.0000 67.2000 ;
	    RECT 125.4000 66.8000 125.8000 67.2000 ;
	    RECT 126.2000 66.8000 126.6000 67.2000 ;
	    RECT 127.0000 67.1000 127.4000 67.2000 ;
	    RECT 127.8000 67.1000 128.1000 67.8000 ;
	    RECT 127.0000 66.8000 128.1000 67.1000 ;
	    RECT 130.2000 67.2000 130.5000 67.8000 ;
	    RECT 130.2000 66.8000 130.6000 67.2000 ;
	    RECT 131.8000 67.1000 132.2000 67.2000 ;
	    RECT 132.6000 67.1000 133.0000 67.2000 ;
	    RECT 131.8000 66.8000 133.0000 67.1000 ;
	    RECT 123.0000 66.2000 123.3000 66.8000 ;
	    RECT 118.2000 65.8000 119.3000 66.1000 ;
	    RECT 119.8000 66.1000 120.2000 66.2000 ;
	    RECT 120.6000 66.1000 121.0000 66.2000 ;
	    RECT 119.8000 65.8000 121.0000 66.1000 ;
	    RECT 123.0000 65.8000 123.4000 66.2000 ;
	    RECT 117.4000 65.2000 117.7000 65.8000 ;
	    RECT 124.6000 65.2000 124.9000 66.8000 ;
	    RECT 133.4000 66.2000 133.7000 67.8000 ;
	    RECT 135.8000 67.2000 136.1000 68.8000 ;
	    RECT 136.6000 67.2000 136.9000 70.8000 ;
	    RECT 135.8000 66.8000 136.2000 67.2000 ;
	    RECT 136.6000 66.8000 137.0000 67.2000 ;
	    RECT 137.4000 66.2000 137.7000 71.8000 ;
	    RECT 138.2000 68.2000 138.5000 74.8000 ;
	    RECT 143.8000 74.2000 144.1000 74.8000 ;
	    RECT 142.2000 73.8000 142.6000 74.2000 ;
	    RECT 143.8000 73.8000 144.2000 74.2000 ;
	    RECT 139.8000 73.1000 140.2000 73.2000 ;
	    RECT 140.6000 73.1000 141.0000 73.2000 ;
	    RECT 139.8000 72.8000 141.0000 73.1000 ;
	    RECT 139.0000 68.8000 139.4000 69.2000 ;
	    RECT 139.0000 68.2000 139.3000 68.8000 ;
	    RECT 138.2000 67.8000 138.6000 68.2000 ;
	    RECT 139.0000 67.8000 139.4000 68.2000 ;
	    RECT 139.8000 67.8000 140.2000 68.2000 ;
	    RECT 139.8000 67.2000 140.1000 67.8000 ;
	    RECT 139.8000 66.8000 140.2000 67.2000 ;
	    RECT 140.6000 66.8000 141.0000 67.2000 ;
	    RECT 140.6000 66.2000 140.9000 66.8000 ;
	    RECT 125.4000 66.1000 125.8000 66.2000 ;
	    RECT 126.2000 66.1000 126.6000 66.2000 ;
	    RECT 125.4000 65.8000 126.6000 66.1000 ;
	    RECT 127.8000 66.1000 128.2000 66.2000 ;
	    RECT 128.6000 66.1000 129.0000 66.2000 ;
	    RECT 127.8000 65.8000 129.0000 66.1000 ;
	    RECT 132.6000 66.1000 133.0000 66.2000 ;
	    RECT 133.4000 66.1000 133.8000 66.2000 ;
	    RECT 132.6000 65.8000 133.8000 66.1000 ;
	    RECT 135.8000 65.8000 136.2000 66.2000 ;
	    RECT 137.4000 66.1000 137.8000 66.2000 ;
	    RECT 138.2000 66.1000 138.6000 66.2000 ;
	    RECT 137.4000 65.8000 138.6000 66.1000 ;
	    RECT 140.6000 65.8000 141.0000 66.2000 ;
	    RECT 141.4000 65.8000 141.8000 66.2000 ;
	    RECT 117.4000 64.8000 117.8000 65.2000 ;
	    RECT 118.2000 65.1000 118.6000 65.2000 ;
	    RECT 119.0000 65.1000 119.4000 65.2000 ;
	    RECT 118.2000 64.8000 119.4000 65.1000 ;
	    RECT 124.6000 64.8000 125.0000 65.2000 ;
	    RECT 129.4000 65.1000 129.8000 65.2000 ;
	    RECT 130.2000 65.1000 130.6000 65.2000 ;
	    RECT 129.4000 64.8000 130.6000 65.1000 ;
	    RECT 133.4000 65.1000 133.8000 65.2000 ;
	    RECT 134.4000 65.1000 134.8000 65.2000 ;
	    RECT 133.4000 64.8000 134.8000 65.1000 ;
	    RECT 111.0000 63.8000 111.4000 64.2000 ;
	    RECT 114.2000 63.8000 114.6000 64.2000 ;
	    RECT 116.6000 63.8000 117.0000 64.2000 ;
	    RECT 120.6000 63.8000 121.0000 64.2000 ;
	    RECT 110.2000 62.8000 110.6000 63.2000 ;
	    RECT 119.8000 62.8000 120.2000 63.2000 ;
	    RECT 119.8000 62.2000 120.1000 62.8000 ;
	    RECT 119.8000 61.8000 120.2000 62.2000 ;
	    RECT 110.2000 60.8000 110.6000 61.2000 ;
	    RECT 110.2000 59.2000 110.5000 60.8000 ;
	    RECT 112.6000 59.8000 113.0000 60.2000 ;
	    RECT 110.2000 58.8000 110.6000 59.2000 ;
	    RECT 108.6000 55.8000 109.7000 56.1000 ;
	    RECT 108.6000 54.8000 109.0000 55.2000 ;
	    RECT 107.8000 52.8000 108.2000 53.2000 ;
	    RECT 108.6000 52.2000 108.9000 54.8000 ;
	    RECT 107.0000 51.8000 107.4000 52.2000 ;
	    RECT 108.6000 51.8000 109.0000 52.2000 ;
	    RECT 104.6000 43.8000 105.0000 44.2000 ;
	    RECT 105.4000 43.1000 105.8000 48.9000 ;
	    RECT 103.0000 41.8000 103.4000 42.2000 ;
	    RECT 103.0000 41.2000 103.3000 41.8000 ;
	    RECT 103.0000 40.8000 103.4000 41.2000 ;
	    RECT 100.6000 37.8000 101.0000 38.2000 ;
	    RECT 105.4000 37.8000 105.8000 38.2000 ;
	    RECT 106.2000 37.8000 106.6000 38.2000 ;
	    RECT 105.4000 36.2000 105.7000 37.8000 ;
	    RECT 102.2000 35.8000 102.6000 36.2000 ;
	    RECT 103.6000 36.1000 104.0000 36.2000 ;
	    RECT 104.6000 36.1000 105.0000 36.2000 ;
	    RECT 103.6000 35.8000 105.0000 36.1000 ;
	    RECT 105.4000 35.8000 105.8000 36.2000 ;
	    RECT 102.2000 34.2000 102.5000 35.8000 ;
	    RECT 106.2000 35.2000 106.5000 37.8000 ;
	    RECT 107.0000 37.2000 107.3000 51.8000 ;
	    RECT 107.8000 46.8000 108.2000 47.2000 ;
	    RECT 107.0000 36.8000 107.4000 37.2000 ;
	    RECT 103.0000 35.1000 103.4000 35.2000 ;
	    RECT 103.8000 35.1000 104.2000 35.2000 ;
	    RECT 103.0000 34.8000 104.2000 35.1000 ;
	    RECT 106.2000 34.8000 106.6000 35.2000 ;
	    RECT 91.8000 33.8000 92.2000 34.2000 ;
	    RECT 94.2000 33.8000 94.6000 34.2000 ;
	    RECT 99.0000 34.1000 99.4000 34.2000 ;
	    RECT 99.8000 34.1000 100.2000 34.2000 ;
	    RECT 99.0000 33.8000 100.2000 34.1000 ;
	    RECT 102.2000 33.8000 102.6000 34.2000 ;
	    RECT 105.4000 33.8000 105.8000 34.2000 ;
	    RECT 91.8000 26.2000 92.1000 33.8000 ;
	    RECT 93.4000 32.8000 93.8000 33.2000 ;
	    RECT 93.4000 29.2000 93.7000 32.8000 ;
	    RECT 93.4000 28.8000 93.8000 29.2000 ;
	    RECT 94.2000 27.2000 94.5000 33.8000 ;
	    RECT 102.2000 33.2000 102.5000 33.8000 ;
	    RECT 105.4000 33.2000 105.7000 33.8000 ;
	    RECT 102.2000 32.8000 102.6000 33.2000 ;
	    RECT 105.4000 32.8000 105.8000 33.2000 ;
	    RECT 94.2000 26.8000 94.6000 27.2000 ;
	    RECT 94.2000 26.2000 94.5000 26.8000 ;
	    RECT 91.8000 25.8000 92.2000 26.2000 ;
	    RECT 94.2000 25.8000 94.6000 26.2000 ;
	    RECT 95.0000 23.1000 95.4000 28.9000 ;
	    RECT 98.2000 28.8000 98.6000 29.2000 ;
	    RECT 96.6000 27.8000 97.0000 28.2000 ;
	    RECT 94.2000 17.8000 94.6000 18.2000 ;
	    RECT 94.2000 15.2000 94.5000 17.8000 ;
	    RECT 96.6000 16.2000 96.9000 27.8000 ;
	    RECT 98.2000 26.2000 98.5000 28.8000 ;
	    RECT 98.2000 25.8000 98.6000 26.2000 ;
	    RECT 102.2000 26.1000 102.6000 26.2000 ;
	    RECT 103.0000 26.1000 103.4000 26.2000 ;
	    RECT 102.2000 25.8000 103.4000 26.1000 ;
	    RECT 104.6000 24.1000 105.0000 24.2000 ;
	    RECT 105.4000 24.1000 105.8000 24.2000 ;
	    RECT 104.6000 23.8000 105.8000 24.1000 ;
	    RECT 107.0000 23.1000 107.4000 28.9000 ;
	    RECT 107.8000 27.2000 108.1000 46.8000 ;
	    RECT 108.6000 45.8000 109.0000 46.2000 ;
	    RECT 108.6000 44.2000 108.9000 45.8000 ;
	    RECT 108.6000 43.8000 109.0000 44.2000 ;
	    RECT 109.4000 39.2000 109.7000 55.8000 ;
	    RECT 111.8000 55.8000 112.2000 56.2000 ;
	    RECT 111.8000 53.2000 112.1000 55.8000 ;
	    RECT 111.8000 52.8000 112.2000 53.2000 ;
	    RECT 110.2000 43.1000 110.6000 48.9000 ;
	    RECT 111.8000 45.1000 112.2000 47.9000 ;
	    RECT 112.6000 47.2000 112.9000 59.8000 ;
	    RECT 119.0000 58.8000 119.4000 59.2000 ;
	    RECT 119.0000 58.2000 119.3000 58.8000 ;
	    RECT 113.4000 57.8000 113.8000 58.2000 ;
	    RECT 119.0000 57.8000 119.4000 58.2000 ;
	    RECT 113.4000 57.2000 113.7000 57.8000 ;
	    RECT 113.4000 56.8000 113.8000 57.2000 ;
	    RECT 119.0000 56.8000 119.4000 57.2000 ;
	    RECT 114.2000 55.8000 114.6000 56.2000 ;
	    RECT 113.4000 54.8000 113.8000 55.2000 ;
	    RECT 113.4000 49.2000 113.7000 54.8000 ;
	    RECT 114.2000 54.2000 114.5000 55.8000 ;
	    RECT 119.0000 55.2000 119.3000 56.8000 ;
	    RECT 115.0000 55.1000 115.4000 55.2000 ;
	    RECT 115.8000 55.1000 116.2000 55.2000 ;
	    RECT 115.0000 54.8000 116.2000 55.1000 ;
	    RECT 119.0000 54.8000 119.4000 55.2000 ;
	    RECT 114.2000 53.8000 114.6000 54.2000 ;
	    RECT 114.2000 51.8000 114.6000 52.2000 ;
	    RECT 113.4000 48.8000 113.8000 49.2000 ;
	    RECT 112.6000 46.8000 113.0000 47.2000 ;
	    RECT 114.2000 46.2000 114.5000 51.8000 ;
	    RECT 114.2000 45.8000 114.6000 46.2000 ;
	    RECT 114.2000 42.1000 114.5000 45.8000 ;
	    RECT 117.4000 45.1000 117.8000 47.9000 ;
	    RECT 118.2000 46.8000 118.6000 47.2000 ;
	    RECT 118.2000 46.2000 118.5000 46.8000 ;
	    RECT 118.2000 45.8000 118.6000 46.2000 ;
	    RECT 119.0000 43.1000 119.4000 48.9000 ;
	    RECT 120.6000 48.2000 120.9000 63.8000 ;
	    RECT 121.4000 58.8000 121.8000 59.2000 ;
	    RECT 121.4000 56.2000 121.7000 58.8000 ;
	    RECT 124.6000 58.2000 124.9000 64.8000 ;
	    RECT 133.4000 63.8000 133.8000 64.2000 ;
	    RECT 130.2000 61.8000 130.6000 62.2000 ;
	    RECT 130.2000 59.2000 130.5000 61.8000 ;
	    RECT 133.4000 59.2000 133.7000 63.8000 ;
	    RECT 130.2000 58.8000 130.6000 59.2000 ;
	    RECT 133.4000 58.8000 133.8000 59.2000 ;
	    RECT 124.6000 57.8000 125.0000 58.2000 ;
	    RECT 125.4000 57.8000 125.8000 58.2000 ;
	    RECT 125.4000 57.2000 125.7000 57.8000 ;
	    RECT 123.0000 56.8000 123.4000 57.2000 ;
	    RECT 125.4000 56.8000 125.8000 57.2000 ;
	    RECT 121.4000 55.8000 121.8000 56.2000 ;
	    RECT 123.0000 54.1000 123.3000 56.8000 ;
	    RECT 123.8000 55.8000 124.2000 56.2000 ;
	    RECT 130.2000 55.8000 130.6000 56.2000 ;
	    RECT 123.8000 55.2000 124.1000 55.8000 ;
	    RECT 130.2000 55.2000 130.5000 55.8000 ;
	    RECT 135.8000 55.2000 136.1000 65.8000 ;
	    RECT 139.0000 65.1000 139.4000 65.2000 ;
	    RECT 139.8000 65.1000 140.2000 65.2000 ;
	    RECT 139.0000 64.8000 140.2000 65.1000 ;
	    RECT 140.6000 55.2000 140.9000 65.8000 ;
	    RECT 141.4000 65.2000 141.7000 65.8000 ;
	    RECT 141.4000 64.8000 141.8000 65.2000 ;
	    RECT 142.2000 64.1000 142.5000 73.8000 ;
	    RECT 145.4000 66.2000 145.7000 76.8000 ;
	    RECT 145.4000 65.8000 145.8000 66.2000 ;
	    RECT 142.2000 63.8000 143.3000 64.1000 ;
	    RECT 123.8000 54.8000 124.2000 55.2000 ;
	    RECT 124.6000 54.8000 125.0000 55.2000 ;
	    RECT 125.4000 54.8000 125.8000 55.2000 ;
	    RECT 127.8000 54.8000 128.2000 55.2000 ;
	    RECT 130.2000 54.8000 130.6000 55.2000 ;
	    RECT 135.8000 54.8000 136.2000 55.2000 ;
	    RECT 137.4000 54.8000 137.8000 55.2000 ;
	    RECT 138.2000 54.8000 138.6000 55.2000 ;
	    RECT 140.6000 54.8000 141.0000 55.2000 ;
	    RECT 142.2000 54.8000 142.6000 55.2000 ;
	    RECT 124.6000 54.2000 124.9000 54.8000 ;
	    RECT 125.4000 54.2000 125.7000 54.8000 ;
	    RECT 127.8000 54.2000 128.1000 54.8000 ;
	    RECT 123.8000 54.1000 124.2000 54.2000 ;
	    RECT 123.0000 53.8000 124.2000 54.1000 ;
	    RECT 124.6000 53.8000 125.0000 54.2000 ;
	    RECT 125.4000 53.8000 125.8000 54.2000 ;
	    RECT 127.0000 54.1000 127.4000 54.2000 ;
	    RECT 127.8000 54.1000 128.2000 54.2000 ;
	    RECT 127.0000 53.8000 128.2000 54.1000 ;
	    RECT 120.6000 47.8000 121.0000 48.2000 ;
	    RECT 114.2000 41.8000 115.3000 42.1000 ;
	    RECT 109.4000 38.8000 109.8000 39.2000 ;
	    RECT 111.0000 36.8000 111.4000 37.2000 ;
	    RECT 111.0000 36.2000 111.3000 36.8000 ;
	    RECT 109.4000 35.8000 109.8000 36.2000 ;
	    RECT 110.2000 35.8000 110.6000 36.2000 ;
	    RECT 111.0000 35.8000 111.4000 36.2000 ;
	    RECT 109.4000 35.2000 109.7000 35.8000 ;
	    RECT 110.2000 35.2000 110.5000 35.8000 ;
	    RECT 109.4000 34.8000 109.8000 35.2000 ;
	    RECT 110.2000 34.8000 110.6000 35.2000 ;
	    RECT 111.8000 33.1000 112.2000 35.9000 ;
	    RECT 112.6000 34.8000 113.0000 35.2000 ;
	    RECT 112.6000 34.2000 112.9000 34.8000 ;
	    RECT 112.6000 33.8000 113.0000 34.2000 ;
	    RECT 113.4000 32.1000 113.8000 37.9000 ;
	    RECT 114.2000 35.8000 114.6000 36.2000 ;
	    RECT 114.2000 35.1000 114.5000 35.8000 ;
	    RECT 114.2000 34.7000 114.6000 35.1000 ;
	    RECT 107.8000 26.8000 108.2000 27.2000 ;
	    RECT 107.8000 26.2000 108.1000 26.8000 ;
	    RECT 107.8000 25.8000 108.2000 26.2000 ;
	    RECT 110.2000 26.1000 110.6000 26.2000 ;
	    RECT 111.0000 26.1000 111.4000 26.3000 ;
	    RECT 110.2000 25.9000 111.4000 26.1000 ;
	    RECT 110.2000 25.8000 111.3000 25.9000 ;
	    RECT 111.8000 23.1000 112.2000 28.9000 ;
	    RECT 113.4000 25.1000 113.8000 27.9000 ;
	    RECT 114.2000 27.8000 114.6000 28.2000 ;
	    RECT 114.2000 24.2000 114.5000 27.8000 ;
	    RECT 114.2000 23.8000 114.6000 24.2000 ;
	    RECT 96.6000 15.8000 97.0000 16.2000 ;
	    RECT 100.6000 15.8000 101.0000 16.2000 ;
	    RECT 111.0000 15.8000 111.4000 16.2000 ;
	    RECT 100.6000 15.2000 100.9000 15.8000 ;
	    RECT 111.0000 15.2000 111.3000 15.8000 ;
	    RECT 91.0000 14.8000 91.4000 15.2000 ;
	    RECT 94.2000 14.8000 94.6000 15.2000 ;
	    RECT 100.6000 14.8000 101.0000 15.2000 ;
	    RECT 101.4000 14.8000 101.8000 15.2000 ;
	    RECT 105.4000 15.1000 105.8000 15.2000 ;
	    RECT 106.2000 15.1000 106.6000 15.2000 ;
	    RECT 105.4000 14.8000 106.6000 15.1000 ;
	    RECT 107.8000 15.1000 108.2000 15.2000 ;
	    RECT 108.6000 15.1000 109.0000 15.2000 ;
	    RECT 107.8000 14.8000 109.0000 15.1000 ;
	    RECT 110.2000 14.8000 110.6000 15.2000 ;
	    RECT 111.0000 14.8000 111.4000 15.2000 ;
	    RECT 101.4000 14.2000 101.7000 14.8000 ;
	    RECT 110.2000 14.2000 110.5000 14.8000 ;
	    RECT 89.4000 13.8000 89.8000 14.2000 ;
	    RECT 95.8000 13.8000 96.2000 14.2000 ;
	    RECT 97.4000 14.1000 97.8000 14.2000 ;
	    RECT 98.2000 14.1000 98.6000 14.2000 ;
	    RECT 97.4000 13.8000 98.6000 14.1000 ;
	    RECT 101.4000 13.8000 101.8000 14.2000 ;
	    RECT 108.6000 13.8000 109.0000 14.2000 ;
	    RECT 110.2000 13.8000 110.6000 14.2000 ;
	    RECT 95.8000 13.2000 96.1000 13.8000 ;
	    RECT 85.4000 12.8000 85.8000 13.2000 ;
	    RECT 93.4000 13.1000 93.8000 13.2000 ;
	    RECT 94.2000 13.1000 94.6000 13.2000 ;
	    RECT 93.4000 12.8000 94.6000 13.1000 ;
	    RECT 95.8000 12.8000 96.2000 13.2000 ;
	    RECT 102.2000 12.8000 102.6000 13.2000 ;
	    RECT 103.8000 12.8000 104.2000 13.2000 ;
	    RECT 106.2000 12.8000 106.6000 13.2000 ;
	    RECT 102.2000 12.2000 102.5000 12.8000 ;
	    RECT 80.6000 11.8000 81.0000 12.2000 ;
	    RECT 86.2000 12.1000 86.6000 12.2000 ;
	    RECT 87.0000 12.1000 87.4000 12.2000 ;
	    RECT 86.2000 11.8000 87.4000 12.1000 ;
	    RECT 87.8000 11.8000 88.2000 12.2000 ;
	    RECT 92.6000 11.8000 93.0000 12.2000 ;
	    RECT 95.0000 11.8000 95.4000 12.2000 ;
	    RECT 102.2000 11.8000 102.6000 12.2000 ;
	    RECT 75.0000 6.1000 75.4000 6.2000 ;
	    RECT 75.8000 6.1000 76.2000 6.2000 ;
	    RECT 75.0000 5.8000 76.2000 6.1000 ;
	    RECT 74.2000 3.8000 74.6000 4.2000 ;
	    RECT 77.4000 3.1000 77.8000 8.9000 ;
	    RECT 79.8000 8.8000 80.2000 9.2000 ;
	    RECT 80.6000 8.2000 80.9000 11.8000 ;
	    RECT 83.8000 9.8000 84.2000 10.2000 ;
	    RECT 78.2000 6.8000 78.6000 7.2000 ;
	    RECT 78.2000 6.2000 78.5000 6.8000 ;
	    RECT 78.2000 5.8000 78.6000 6.2000 ;
	    RECT 79.0000 5.1000 79.4000 7.9000 ;
	    RECT 80.6000 7.8000 81.0000 8.2000 ;
	    RECT 81.4000 7.8000 81.8000 8.2000 ;
	    RECT 81.4000 6.2000 81.7000 7.8000 ;
	    RECT 83.8000 6.2000 84.1000 9.8000 ;
	    RECT 81.4000 5.8000 81.8000 6.2000 ;
	    RECT 83.8000 5.8000 84.2000 6.2000 ;
	    RECT 84.6000 5.1000 85.0000 7.9000 ;
	    RECT 86.2000 3.1000 86.6000 8.9000 ;
	    RECT 87.8000 6.2000 88.1000 11.8000 ;
	    RECT 90.2000 6.8000 90.6000 7.2000 ;
	    RECT 90.2000 6.2000 90.5000 6.8000 ;
	    RECT 87.8000 5.8000 88.2000 6.2000 ;
	    RECT 90.2000 5.8000 90.6000 6.2000 ;
	    RECT 91.0000 3.1000 91.4000 8.9000 ;
	    RECT 92.6000 8.2000 92.9000 11.8000 ;
	    RECT 95.0000 10.2000 95.3000 11.8000 ;
	    RECT 95.0000 9.8000 95.4000 10.2000 ;
	    RECT 103.8000 9.2000 104.1000 12.8000 ;
	    RECT 93.4000 8.8000 93.8000 9.2000 ;
	    RECT 93.4000 8.2000 93.7000 8.8000 ;
	    RECT 92.6000 7.8000 93.0000 8.2000 ;
	    RECT 93.4000 7.8000 93.8000 8.2000 ;
	    RECT 96.6000 5.8000 97.0000 6.2000 ;
	    RECT 96.6000 4.2000 96.9000 5.8000 ;
	    RECT 96.6000 3.8000 97.0000 4.2000 ;
	    RECT 99.8000 4.1000 100.2000 4.2000 ;
	    RECT 100.6000 4.1000 101.0000 4.2000 ;
	    RECT 99.8000 3.8000 101.0000 4.1000 ;
	    RECT 103.0000 3.1000 103.4000 8.9000 ;
	    RECT 103.8000 8.8000 104.2000 9.2000 ;
	    RECT 103.8000 6.1000 104.2000 6.2000 ;
	    RECT 104.6000 6.1000 105.0000 6.2000 ;
	    RECT 103.8000 5.8000 105.0000 6.1000 ;
	    RECT 106.2000 4.2000 106.5000 12.8000 ;
	    RECT 107.0000 10.8000 107.4000 11.2000 ;
	    RECT 107.0000 8.2000 107.3000 10.8000 ;
	    RECT 107.0000 7.8000 107.4000 8.2000 ;
	    RECT 107.0000 6.8000 107.4000 7.2000 ;
	    RECT 107.0000 6.3000 107.3000 6.8000 ;
	    RECT 107.0000 5.9000 107.4000 6.3000 ;
	    RECT 107.0000 5.8000 107.3000 5.9000 ;
	    RECT 106.2000 3.8000 106.6000 4.2000 ;
	    RECT 107.8000 3.1000 108.2000 8.9000 ;
	    RECT 108.6000 6.2000 108.9000 13.8000 ;
	    RECT 114.2000 13.2000 114.5000 23.8000 ;
	    RECT 115.0000 15.2000 115.3000 41.8000 ;
	    RECT 115.8000 41.8000 116.2000 42.2000 ;
	    RECT 115.8000 36.2000 116.1000 41.8000 ;
	    RECT 120.6000 39.2000 120.9000 47.8000 ;
	    RECT 121.4000 46.8000 121.8000 47.2000 ;
	    RECT 121.4000 46.2000 121.7000 46.8000 ;
	    RECT 121.4000 45.8000 121.8000 46.2000 ;
	    RECT 123.8000 43.1000 124.2000 48.9000 ;
	    RECT 124.6000 46.2000 124.9000 53.8000 ;
	    RECT 130.2000 51.2000 130.5000 54.8000 ;
	    RECT 131.0000 54.1000 131.4000 54.2000 ;
	    RECT 131.8000 54.1000 132.2000 54.2000 ;
	    RECT 131.0000 53.8000 132.2000 54.1000 ;
	    RECT 131.8000 53.1000 132.2000 53.2000 ;
	    RECT 132.6000 53.1000 133.0000 53.2000 ;
	    RECT 131.8000 52.8000 133.0000 53.1000 ;
	    RECT 131.8000 51.8000 132.2000 52.2000 ;
	    RECT 130.2000 50.8000 130.6000 51.2000 ;
	    RECT 126.2000 49.1000 126.6000 49.2000 ;
	    RECT 127.0000 49.1000 127.4000 49.2000 ;
	    RECT 126.2000 48.8000 127.4000 49.1000 ;
	    RECT 130.2000 48.8000 130.6000 49.2000 ;
	    RECT 130.2000 48.2000 130.5000 48.8000 ;
	    RECT 130.2000 47.8000 130.6000 48.2000 ;
	    RECT 127.8000 46.8000 128.2000 47.2000 ;
	    RECT 128.6000 47.1000 129.0000 47.2000 ;
	    RECT 129.4000 47.1000 129.8000 47.2000 ;
	    RECT 128.6000 46.8000 129.8000 47.1000 ;
	    RECT 131.8000 47.1000 132.1000 51.8000 ;
	    RECT 135.8000 51.2000 136.1000 54.8000 ;
	    RECT 137.4000 54.1000 137.7000 54.8000 ;
	    RECT 136.6000 53.8000 137.7000 54.1000 ;
	    RECT 134.2000 50.8000 134.6000 51.2000 ;
	    RECT 135.8000 50.8000 136.2000 51.2000 ;
	    RECT 133.4000 49.8000 133.8000 50.2000 ;
	    RECT 131.8000 46.8000 132.9000 47.1000 ;
	    RECT 127.8000 46.2000 128.1000 46.8000 ;
	    RECT 124.6000 45.8000 125.0000 46.2000 ;
	    RECT 126.2000 46.1000 126.6000 46.2000 ;
	    RECT 127.0000 46.1000 127.4000 46.2000 ;
	    RECT 126.2000 45.8000 127.4000 46.1000 ;
	    RECT 127.8000 45.8000 128.2000 46.2000 ;
	    RECT 131.0000 46.1000 131.4000 46.2000 ;
	    RECT 131.8000 46.1000 132.2000 46.2000 ;
	    RECT 131.0000 45.8000 132.2000 46.1000 ;
	    RECT 120.6000 38.8000 121.0000 39.2000 ;
	    RECT 121.4000 38.8000 121.8000 39.2000 ;
	    RECT 120.6000 38.2000 120.9000 38.8000 ;
	    RECT 115.8000 35.8000 116.2000 36.2000 ;
	    RECT 118.2000 32.1000 118.6000 37.9000 ;
	    RECT 120.6000 37.8000 121.0000 38.2000 ;
	    RECT 121.4000 35.2000 121.7000 38.8000 ;
	    RECT 122.2000 35.8000 122.6000 36.2000 ;
	    RECT 121.4000 34.8000 121.8000 35.2000 ;
	    RECT 122.2000 34.2000 122.5000 35.8000 ;
	    RECT 122.2000 33.8000 122.6000 34.2000 ;
	    RECT 123.8000 32.8000 124.2000 33.2000 ;
	    RECT 124.6000 33.1000 125.0000 35.9000 ;
	    RECT 125.4000 34.8000 125.8000 35.2000 ;
	    RECT 125.4000 34.2000 125.7000 34.8000 ;
	    RECT 125.4000 33.8000 125.8000 34.2000 ;
	    RECT 123.8000 32.2000 124.1000 32.8000 ;
	    RECT 123.0000 31.8000 123.4000 32.2000 ;
	    RECT 123.8000 31.8000 124.2000 32.2000 ;
	    RECT 126.2000 32.1000 126.6000 37.9000 ;
	    RECT 127.8000 36.2000 128.1000 45.8000 ;
	    RECT 132.6000 45.2000 132.9000 46.8000 ;
	    RECT 132.6000 44.8000 133.0000 45.2000 ;
	    RECT 133.4000 39.2000 133.7000 49.8000 ;
	    RECT 134.2000 46.2000 134.5000 50.8000 ;
	    RECT 135.8000 48.1000 136.2000 48.2000 ;
	    RECT 136.6000 48.1000 136.9000 53.8000 ;
	    RECT 135.8000 47.8000 136.9000 48.1000 ;
	    RECT 135.0000 47.1000 135.4000 47.2000 ;
	    RECT 135.8000 47.1000 136.2000 47.2000 ;
	    RECT 135.0000 46.8000 136.2000 47.1000 ;
	    RECT 138.2000 46.2000 138.5000 54.8000 ;
	    RECT 140.6000 54.2000 140.9000 54.8000 ;
	    RECT 140.6000 53.8000 141.0000 54.2000 ;
	    RECT 141.4000 51.8000 141.8000 52.2000 ;
	    RECT 140.6000 48.8000 141.0000 49.2000 ;
	    RECT 139.0000 47.1000 139.4000 47.2000 ;
	    RECT 139.8000 47.1000 140.2000 47.2000 ;
	    RECT 139.0000 46.8000 140.2000 47.1000 ;
	    RECT 140.6000 46.2000 140.9000 48.8000 ;
	    RECT 134.2000 45.8000 134.6000 46.2000 ;
	    RECT 138.2000 45.8000 138.6000 46.2000 ;
	    RECT 140.6000 45.8000 141.0000 46.2000 ;
	    RECT 141.4000 45.2000 141.7000 51.8000 ;
	    RECT 142.2000 50.2000 142.5000 54.8000 ;
	    RECT 143.0000 53.2000 143.3000 63.8000 ;
	    RECT 143.8000 61.8000 144.2000 62.2000 ;
	    RECT 143.8000 54.2000 144.1000 61.8000 ;
	    RECT 146.2000 59.2000 146.5000 103.8000 ;
	    RECT 146.2000 58.8000 146.6000 59.2000 ;
	    RECT 145.4000 54.8000 145.8000 55.2000 ;
	    RECT 145.4000 54.2000 145.7000 54.8000 ;
	    RECT 143.8000 53.8000 144.2000 54.2000 ;
	    RECT 145.4000 53.8000 145.8000 54.2000 ;
	    RECT 143.0000 52.8000 143.4000 53.2000 ;
	    RECT 145.4000 52.8000 145.8000 53.2000 ;
	    RECT 142.2000 49.8000 142.6000 50.2000 ;
	    RECT 145.4000 49.2000 145.7000 52.8000 ;
	    RECT 145.4000 48.8000 145.8000 49.2000 ;
	    RECT 144.6000 46.1000 145.0000 46.2000 ;
	    RECT 143.8000 45.8000 145.0000 46.1000 ;
	    RECT 139.8000 45.1000 140.2000 45.2000 ;
	    RECT 140.6000 45.1000 141.0000 45.2000 ;
	    RECT 139.8000 44.8000 141.0000 45.1000 ;
	    RECT 141.4000 44.8000 141.8000 45.2000 ;
	    RECT 139.8000 43.8000 140.2000 44.2000 ;
	    RECT 134.2000 41.8000 134.6000 42.2000 ;
	    RECT 136.6000 41.8000 137.0000 42.2000 ;
	    RECT 133.4000 38.8000 133.8000 39.2000 ;
	    RECT 127.8000 35.8000 128.2000 36.2000 ;
	    RECT 127.8000 35.1000 128.2000 35.2000 ;
	    RECT 128.6000 35.1000 129.0000 35.2000 ;
	    RECT 127.8000 34.8000 129.0000 35.1000 ;
	    RECT 128.6000 32.8000 129.0000 33.2000 ;
	    RECT 115.8000 26.8000 116.2000 27.2000 ;
	    RECT 115.8000 26.2000 116.1000 26.8000 ;
	    RECT 115.8000 25.8000 116.2000 26.2000 ;
	    RECT 117.4000 25.8000 117.8000 26.2000 ;
	    RECT 115.0000 14.8000 115.4000 15.2000 ;
	    RECT 117.4000 14.2000 117.7000 25.8000 ;
	    RECT 118.2000 25.1000 118.6000 27.9000 ;
	    RECT 119.0000 27.8000 119.4000 28.2000 ;
	    RECT 119.0000 27.2000 119.3000 27.8000 ;
	    RECT 119.0000 26.8000 119.4000 27.2000 ;
	    RECT 119.8000 23.1000 120.2000 28.9000 ;
	    RECT 123.0000 26.2000 123.3000 31.8000 ;
	    RECT 128.6000 29.2000 128.9000 32.8000 ;
	    RECT 131.0000 32.1000 131.4000 37.9000 ;
	    RECT 134.2000 37.2000 134.5000 41.8000 ;
	    RECT 134.2000 36.8000 134.6000 37.2000 ;
	    RECT 135.0000 35.8000 135.4000 36.2000 ;
	    RECT 131.8000 34.8000 132.2000 35.2000 ;
	    RECT 133.4000 35.1000 133.8000 35.2000 ;
	    RECT 134.2000 35.1000 134.6000 35.2000 ;
	    RECT 133.4000 34.8000 134.6000 35.1000 ;
	    RECT 131.8000 29.2000 132.1000 34.8000 ;
	    RECT 135.0000 34.2000 135.3000 35.8000 ;
	    RECT 136.6000 35.2000 136.9000 41.8000 ;
	    RECT 139.8000 39.2000 140.1000 43.8000 ;
	    RECT 139.8000 38.8000 140.2000 39.2000 ;
	    RECT 137.4000 35.8000 137.8000 36.2000 ;
	    RECT 137.4000 35.2000 137.7000 35.8000 ;
	    RECT 143.8000 35.2000 144.1000 45.8000 ;
	    RECT 136.6000 34.8000 137.0000 35.2000 ;
	    RECT 137.4000 34.8000 137.8000 35.2000 ;
	    RECT 141.4000 34.8000 141.8000 35.2000 ;
	    RECT 143.8000 34.8000 144.2000 35.2000 ;
	    RECT 135.0000 33.8000 135.4000 34.2000 ;
	    RECT 136.6000 33.8000 137.0000 34.2000 ;
	    RECT 140.6000 33.8000 141.0000 34.2000 ;
	    RECT 133.4000 31.8000 133.8000 32.2000 ;
	    RECT 135.8000 31.8000 136.2000 32.2000 ;
	    RECT 133.4000 29.2000 133.7000 31.8000 ;
	    RECT 135.8000 29.2000 136.1000 31.8000 ;
	    RECT 123.0000 25.8000 123.4000 26.2000 ;
	    RECT 124.6000 23.1000 125.0000 28.9000 ;
	    RECT 127.0000 28.8000 127.4000 29.2000 ;
	    RECT 128.6000 28.8000 129.0000 29.2000 ;
	    RECT 131.8000 28.8000 132.2000 29.2000 ;
	    RECT 133.4000 28.8000 133.8000 29.2000 ;
	    RECT 135.0000 28.8000 135.4000 29.2000 ;
	    RECT 135.8000 28.8000 136.2000 29.2000 ;
	    RECT 127.0000 28.2000 127.3000 28.8000 ;
	    RECT 135.0000 28.2000 135.3000 28.8000 ;
	    RECT 127.0000 27.8000 127.4000 28.2000 ;
	    RECT 129.4000 28.1000 129.8000 28.2000 ;
	    RECT 130.2000 28.1000 130.6000 28.2000 ;
	    RECT 129.4000 27.8000 130.6000 28.1000 ;
	    RECT 135.0000 27.8000 135.4000 28.2000 ;
	    RECT 130.2000 26.8000 130.6000 27.2000 ;
	    RECT 131.0000 26.8000 131.4000 27.2000 ;
	    RECT 130.2000 26.2000 130.5000 26.8000 ;
	    RECT 131.0000 26.2000 131.3000 26.8000 ;
	    RECT 127.0000 26.1000 127.4000 26.2000 ;
	    RECT 127.8000 26.1000 128.2000 26.2000 ;
	    RECT 127.0000 25.8000 128.2000 26.1000 ;
	    RECT 130.2000 25.8000 130.6000 26.2000 ;
	    RECT 131.0000 25.8000 131.4000 26.2000 ;
	    RECT 132.6000 26.1000 133.0000 26.2000 ;
	    RECT 133.4000 26.1000 133.8000 26.2000 ;
	    RECT 132.6000 25.8000 133.8000 26.1000 ;
	    RECT 120.6000 16.8000 121.0000 17.2000 ;
	    RECT 124.6000 16.8000 125.0000 17.2000 ;
	    RECT 120.6000 15.2000 120.9000 16.8000 ;
	    RECT 121.4000 15.8000 121.8000 16.2000 ;
	    RECT 121.4000 15.2000 121.7000 15.8000 ;
	    RECT 120.6000 14.8000 121.0000 15.2000 ;
	    RECT 121.4000 14.8000 121.8000 15.2000 ;
	    RECT 123.0000 14.8000 123.4000 15.2000 ;
	    RECT 123.0000 14.2000 123.3000 14.8000 ;
	    RECT 117.4000 13.8000 117.8000 14.2000 ;
	    RECT 123.0000 13.8000 123.4000 14.2000 ;
	    RECT 124.6000 13.2000 124.9000 16.8000 ;
	    RECT 110.2000 12.8000 110.6000 13.2000 ;
	    RECT 114.2000 12.8000 114.6000 13.2000 ;
	    RECT 124.6000 12.8000 125.0000 13.2000 ;
	    RECT 108.6000 5.8000 109.0000 6.2000 ;
	    RECT 109.4000 5.1000 109.8000 7.9000 ;
	    RECT 110.2000 6.2000 110.5000 12.8000 ;
	    RECT 119.0000 11.8000 119.4000 12.2000 ;
	    RECT 119.0000 10.1000 119.3000 11.8000 ;
	    RECT 119.0000 9.8000 120.1000 10.1000 ;
	    RECT 119.8000 6.2000 120.1000 9.8000 ;
	    RECT 124.6000 6.2000 124.9000 12.8000 ;
	    RECT 127.0000 7.2000 127.3000 25.8000 ;
	    RECT 135.8000 25.1000 136.2000 27.9000 ;
	    RECT 136.6000 27.2000 136.9000 33.8000 ;
	    RECT 140.6000 33.2000 140.9000 33.8000 ;
	    RECT 141.4000 33.2000 141.7000 34.8000 ;
	    RECT 139.0000 33.1000 139.4000 33.2000 ;
	    RECT 139.8000 33.1000 140.2000 33.2000 ;
	    RECT 139.0000 32.8000 140.2000 33.1000 ;
	    RECT 140.6000 32.8000 141.0000 33.2000 ;
	    RECT 141.4000 32.8000 141.8000 33.2000 ;
	    RECT 143.8000 32.2000 144.1000 34.8000 ;
	    RECT 144.6000 32.8000 145.0000 33.2000 ;
	    RECT 143.8000 31.8000 144.2000 32.2000 ;
	    RECT 144.6000 29.2000 144.9000 32.8000 ;
	    RECT 146.2000 31.8000 146.6000 32.2000 ;
	    RECT 136.6000 26.8000 137.0000 27.2000 ;
	    RECT 137.4000 23.1000 137.8000 28.9000 ;
	    RECT 139.0000 28.8000 139.4000 29.2000 ;
	    RECT 138.2000 26.8000 138.6000 27.2000 ;
	    RECT 127.8000 12.1000 128.2000 17.9000 ;
	    RECT 128.6000 15.1000 129.0000 15.2000 ;
	    RECT 129.4000 15.1000 129.8000 15.2000 ;
	    RECT 128.6000 14.8000 129.8000 15.1000 ;
	    RECT 130.2000 14.8000 130.6000 15.2000 ;
	    RECT 130.2000 9.2000 130.5000 14.8000 ;
	    RECT 131.8000 11.8000 132.2000 12.2000 ;
	    RECT 132.6000 12.1000 133.0000 17.9000 ;
	    RECT 134.2000 13.1000 134.6000 15.9000 ;
	    RECT 135.0000 13.1000 135.4000 15.9000 ;
	    RECT 136.6000 12.1000 137.0000 17.9000 ;
	    RECT 137.4000 14.7000 137.8000 15.1000 ;
	    RECT 137.4000 14.2000 137.7000 14.7000 ;
	    RECT 138.2000 14.2000 138.5000 26.8000 ;
	    RECT 139.0000 26.2000 139.3000 28.8000 ;
	    RECT 139.0000 25.8000 139.4000 26.2000 ;
	    RECT 142.2000 23.1000 142.6000 28.9000 ;
	    RECT 144.6000 28.8000 145.0000 29.2000 ;
	    RECT 145.4000 27.8000 145.8000 28.2000 ;
	    RECT 145.4000 26.2000 145.7000 27.8000 ;
	    RECT 145.4000 25.8000 145.8000 26.2000 ;
	    RECT 145.4000 24.8000 145.8000 25.2000 ;
	    RECT 137.4000 13.8000 137.8000 14.2000 ;
	    RECT 138.2000 13.8000 138.6000 14.2000 ;
	    RECT 141.4000 12.1000 141.8000 17.9000 ;
	    RECT 143.8000 15.1000 144.2000 15.2000 ;
	    RECT 144.6000 15.1000 145.0000 15.2000 ;
	    RECT 143.8000 14.8000 145.0000 15.1000 ;
	    RECT 143.0000 12.1000 143.4000 12.2000 ;
	    RECT 143.8000 12.1000 144.2000 12.2000 ;
	    RECT 143.0000 11.8000 144.2000 12.1000 ;
	    RECT 130.2000 8.8000 130.6000 9.2000 ;
	    RECT 127.9000 7.8000 128.3000 7.9000 ;
	    RECT 127.9000 7.5000 130.7000 7.8000 ;
	    RECT 131.0000 7.5000 131.4000 7.9000 ;
	    RECT 127.0000 6.8000 127.4000 7.2000 ;
	    RECT 110.2000 5.8000 110.6000 6.2000 ;
	    RECT 112.6000 6.1000 113.0000 6.2000 ;
	    RECT 113.4000 6.1000 113.8000 6.2000 ;
	    RECT 112.6000 5.8000 113.8000 6.1000 ;
	    RECT 115.0000 6.1000 115.4000 6.2000 ;
	    RECT 115.8000 6.1000 116.2000 6.2000 ;
	    RECT 115.0000 5.8000 116.2000 6.1000 ;
	    RECT 117.4000 6.1000 117.8000 6.2000 ;
	    RECT 118.2000 6.1000 118.6000 6.2000 ;
	    RECT 117.4000 5.8000 118.6000 6.1000 ;
	    RECT 119.8000 5.8000 120.2000 6.2000 ;
	    RECT 121.4000 6.1000 121.8000 6.2000 ;
	    RECT 122.2000 6.1000 122.6000 6.2000 ;
	    RECT 121.4000 5.8000 122.6000 6.1000 ;
	    RECT 124.6000 5.8000 125.0000 6.2000 ;
	    RECT 127.9000 5.1000 128.2000 7.5000 ;
	    RECT 128.6000 7.4000 129.0000 7.5000 ;
	    RECT 130.3000 7.4000 130.7000 7.5000 ;
	    RECT 131.1000 7.1000 131.4000 7.5000 ;
	    RECT 128.6000 6.8000 131.4000 7.1000 ;
	    RECT 131.8000 7.2000 132.1000 11.8000 ;
	    RECT 145.4000 9.2000 145.7000 24.8000 ;
	    RECT 146.2000 19.2000 146.5000 31.8000 ;
	    RECT 146.2000 18.8000 146.6000 19.2000 ;
	    RECT 146.2000 11.8000 146.6000 12.2000 ;
	    RECT 145.4000 8.8000 145.8000 9.2000 ;
	    RECT 144.6000 7.8000 145.0000 8.2000 ;
	    RECT 144.6000 7.2000 144.9000 7.8000 ;
	    RECT 131.8000 6.8000 132.2000 7.2000 ;
	    RECT 144.6000 6.8000 145.0000 7.2000 ;
	    RECT 128.6000 6.1000 128.9000 6.8000 ;
	    RECT 128.5000 5.7000 128.9000 6.1000 ;
	    RECT 131.1000 5.1000 131.4000 6.8000 ;
	    RECT 146.2000 6.2000 146.5000 11.8000 ;
	    RECT 137.4000 6.1000 137.8000 6.2000 ;
	    RECT 138.2000 6.1000 138.6000 6.2000 ;
	    RECT 137.4000 5.8000 138.6000 6.1000 ;
	    RECT 139.8000 6.1000 140.2000 6.2000 ;
	    RECT 140.6000 6.1000 141.0000 6.2000 ;
	    RECT 139.8000 5.8000 141.0000 6.1000 ;
	    RECT 142.2000 6.1000 142.6000 6.2000 ;
	    RECT 143.0000 6.1000 143.4000 6.2000 ;
	    RECT 142.2000 5.8000 143.4000 6.1000 ;
	    RECT 146.2000 5.8000 146.6000 6.2000 ;
	    RECT 127.9000 4.7000 128.3000 5.1000 ;
	    RECT 131.0000 4.7000 131.4000 5.1000 ;
         LAYER metal3 ;
	    RECT 19.8000 117.1000 20.2000 117.2000 ;
	    RECT 21.4000 117.1000 21.8000 117.2000 ;
	    RECT 31.8000 117.1000 32.2000 117.2000 ;
	    RECT 19.8000 116.8000 32.2000 117.1000 ;
	    RECT 7.0000 115.8000 7.4000 116.2000 ;
	    RECT 14.2000 115.8000 14.6000 116.2000 ;
	    RECT 40.6000 116.1000 41.0000 116.2000 ;
	    RECT 42.2000 116.1000 42.6000 116.2000 ;
	    RECT 40.6000 115.8000 42.6000 116.1000 ;
	    RECT 63.8000 115.8000 64.2000 116.2000 ;
	    RECT 65.4000 116.1000 65.8000 116.2000 ;
	    RECT 66.2000 116.1000 66.6000 116.2000 ;
	    RECT 65.4000 115.8000 66.6000 116.1000 ;
	    RECT 73.4000 115.8000 73.8000 116.2000 ;
	    RECT 7.0000 115.1000 7.3000 115.8000 ;
	    RECT 14.2000 115.1000 14.5000 115.8000 ;
	    RECT 7.0000 114.8000 14.5000 115.1000 ;
	    RECT 17.4000 115.1000 17.8000 115.2000 ;
	    RECT 39.0000 115.1000 39.4000 115.2000 ;
	    RECT 17.4000 114.8000 39.4000 115.1000 ;
	    RECT 41.4000 114.8000 41.8000 115.2000 ;
	    RECT 43.8000 115.1000 44.2000 115.2000 ;
	    RECT 52.6000 115.1000 53.0000 115.2000 ;
	    RECT 43.8000 114.8000 53.0000 115.1000 ;
	    RECT 63.8000 115.1000 64.1000 115.8000 ;
	    RECT 73.4000 115.1000 73.7000 115.8000 ;
	    RECT 63.8000 114.8000 73.7000 115.1000 ;
	    RECT 85.4000 115.1000 85.8000 115.2000 ;
	    RECT 87.0000 115.1000 87.4000 115.2000 ;
	    RECT 89.4000 115.1000 89.8000 115.2000 ;
	    RECT 85.4000 114.8000 89.8000 115.1000 ;
	    RECT 117.4000 115.1000 117.8000 115.2000 ;
	    RECT 141.4000 115.1000 141.8000 115.2000 ;
	    RECT 143.8000 115.1000 144.2000 115.2000 ;
	    RECT 144.6000 115.1000 145.0000 115.2000 ;
	    RECT 117.4000 114.8000 129.7000 115.1000 ;
	    RECT 141.4000 114.8000 145.0000 115.1000 ;
	    RECT 38.2000 114.1000 38.6000 114.2000 ;
	    RECT 41.4000 114.1000 41.7000 114.8000 ;
	    RECT 129.4000 114.2000 129.7000 114.8000 ;
	    RECT 38.2000 113.8000 41.7000 114.1000 ;
	    RECT 45.4000 113.8000 45.8000 114.2000 ;
	    RECT 79.0000 114.1000 79.4000 114.2000 ;
	    RECT 67.8000 113.8000 79.4000 114.1000 ;
	    RECT 107.8000 114.1000 108.2000 114.2000 ;
	    RECT 109.4000 114.1000 109.8000 114.2000 ;
	    RECT 107.8000 113.8000 109.8000 114.1000 ;
	    RECT 115.0000 114.1000 115.4000 114.2000 ;
	    RECT 123.8000 114.1000 124.2000 114.2000 ;
	    RECT 115.0000 113.8000 124.2000 114.1000 ;
	    RECT 129.4000 114.1000 129.8000 114.2000 ;
	    RECT 139.8000 114.1000 140.2000 114.2000 ;
	    RECT 129.4000 113.8000 140.2000 114.1000 ;
	    RECT 0.6000 113.1000 1.0000 113.2000 ;
	    RECT 12.6000 113.1000 13.0000 113.2000 ;
	    RECT 17.4000 113.1000 17.8000 113.2000 ;
	    RECT 0.6000 112.8000 17.8000 113.1000 ;
	    RECT 19.0000 112.8000 19.4000 113.2000 ;
	    RECT 36.6000 113.1000 37.0000 113.2000 ;
	    RECT 44.6000 113.1000 45.0000 113.2000 ;
	    RECT 36.6000 112.8000 45.0000 113.1000 ;
	    RECT 45.4000 113.1000 45.7000 113.8000 ;
	    RECT 67.8000 113.2000 68.1000 113.8000 ;
	    RECT 55.8000 113.1000 56.2000 113.2000 ;
	    RECT 45.4000 112.8000 56.2000 113.1000 ;
	    RECT 67.0000 113.1000 67.4000 113.2000 ;
	    RECT 67.8000 113.1000 68.2000 113.2000 ;
	    RECT 67.0000 112.8000 68.2000 113.1000 ;
	    RECT 19.0000 112.1000 19.3000 112.8000 ;
	    RECT 40.6000 112.1000 41.0000 112.2000 ;
	    RECT 51.8000 112.1000 52.2000 112.2000 ;
	    RECT 19.0000 111.8000 52.2000 112.1000 ;
	    RECT 55.0000 112.1000 55.4000 112.2000 ;
	    RECT 58.2000 112.1000 58.6000 112.2000 ;
	    RECT 59.8000 112.1000 60.2000 112.2000 ;
	    RECT 55.0000 111.8000 60.2000 112.1000 ;
	    RECT 97.4000 112.1000 97.8000 112.2000 ;
	    RECT 101.4000 112.1000 101.8000 112.2000 ;
	    RECT 97.4000 111.8000 101.8000 112.1000 ;
	    RECT 28.6000 111.1000 29.0000 111.2000 ;
	    RECT 33.4000 111.1000 33.8000 111.2000 ;
	    RECT 28.6000 110.8000 33.8000 111.1000 ;
	    RECT 37.4000 111.1000 37.8000 111.2000 ;
	    RECT 43.0000 111.1000 43.4000 111.2000 ;
	    RECT 37.4000 110.8000 43.4000 111.1000 ;
	    RECT 54.2000 111.1000 54.6000 111.2000 ;
	    RECT 63.0000 111.1000 63.4000 111.2000 ;
	    RECT 54.2000 110.8000 63.4000 111.1000 ;
	    RECT 75.0000 111.1000 75.4000 111.2000 ;
	    RECT 78.2000 111.1000 78.6000 111.2000 ;
	    RECT 87.8000 111.1000 88.2000 111.2000 ;
	    RECT 75.0000 110.8000 88.2000 111.1000 ;
	    RECT 104.6000 111.1000 105.0000 111.2000 ;
	    RECT 106.2000 111.1000 106.6000 111.2000 ;
	    RECT 104.6000 110.8000 106.6000 111.1000 ;
	    RECT 108.6000 111.1000 109.0000 111.2000 ;
	    RECT 114.2000 111.1000 114.6000 111.2000 ;
	    RECT 108.6000 110.8000 114.6000 111.1000 ;
	    RECT 102.2000 110.1000 102.6000 110.2000 ;
	    RECT 107.0000 110.1000 107.4000 110.2000 ;
	    RECT 102.2000 109.8000 107.4000 110.1000 ;
	    RECT 109.4000 110.1000 109.8000 110.2000 ;
	    RECT 113.4000 110.1000 113.8000 110.2000 ;
	    RECT 109.4000 109.8000 113.8000 110.1000 ;
	    RECT 67.8000 109.1000 68.2000 109.2000 ;
	    RECT 68.6000 109.1000 69.0000 109.2000 ;
	    RECT 74.2000 109.1000 74.6000 109.2000 ;
	    RECT 67.8000 108.8000 74.6000 109.1000 ;
	    RECT 88.6000 109.1000 89.0000 109.2000 ;
	    RECT 92.6000 109.1000 93.0000 109.2000 ;
	    RECT 95.0000 109.1000 95.4000 109.2000 ;
	    RECT 107.8000 109.1000 108.2000 109.2000 ;
	    RECT 88.6000 108.8000 108.2000 109.1000 ;
	    RECT 108.6000 108.8000 109.0000 109.2000 ;
	    RECT 129.4000 109.1000 129.8000 109.2000 ;
	    RECT 134.2000 109.1000 134.6000 109.2000 ;
	    RECT 129.4000 108.8000 134.6000 109.1000 ;
	    RECT 135.8000 109.1000 136.2000 109.2000 ;
	    RECT 140.6000 109.1000 141.0000 109.2000 ;
	    RECT 147.0000 109.1000 147.4000 109.2000 ;
	    RECT 135.8000 108.8000 147.4000 109.1000 ;
	    RECT 6.2000 107.8000 12.9000 108.1000 ;
	    RECT 6.2000 107.2000 6.5000 107.8000 ;
	    RECT 12.6000 107.2000 12.9000 107.8000 ;
	    RECT 28.6000 107.8000 29.0000 108.2000 ;
	    RECT 39.8000 108.1000 40.2000 108.2000 ;
	    RECT 46.2000 108.1000 46.6000 108.2000 ;
	    RECT 39.8000 107.8000 46.6000 108.1000 ;
	    RECT 52.6000 108.1000 53.0000 108.2000 ;
	    RECT 67.0000 108.1000 67.4000 108.2000 ;
	    RECT 52.6000 107.8000 67.4000 108.1000 ;
	    RECT 108.6000 108.1000 108.9000 108.8000 ;
	    RECT 116.6000 108.1000 117.0000 108.2000 ;
	    RECT 108.6000 107.8000 117.0000 108.1000 ;
	    RECT 120.6000 108.1000 121.0000 108.2000 ;
	    RECT 124.6000 108.1000 125.0000 108.2000 ;
	    RECT 139.0000 108.1000 139.4000 108.2000 ;
	    RECT 120.6000 107.8000 125.0000 108.1000 ;
	    RECT 138.2000 107.8000 139.4000 108.1000 ;
	    RECT 6.2000 106.8000 6.6000 107.2000 ;
	    RECT 12.6000 106.8000 13.0000 107.2000 ;
	    RECT 19.8000 107.1000 20.2000 107.2000 ;
	    RECT 28.6000 107.1000 28.9000 107.8000 ;
	    RECT 138.2000 107.2000 138.5000 107.8000 ;
	    RECT 37.4000 107.1000 37.8000 107.2000 ;
	    RECT 47.0000 107.1000 47.4000 107.2000 ;
	    RECT 51.0000 107.1000 51.4000 107.2000 ;
	    RECT 19.8000 106.8000 37.8000 107.1000 ;
	    RECT 41.4000 106.8000 51.4000 107.1000 ;
	    RECT 55.8000 107.1000 56.2000 107.2000 ;
	    RECT 58.2000 107.1000 58.6000 107.2000 ;
	    RECT 61.4000 107.1000 61.8000 107.2000 ;
	    RECT 55.8000 106.8000 61.8000 107.1000 ;
	    RECT 92.6000 107.1000 93.0000 107.2000 ;
	    RECT 105.4000 107.1000 105.8000 107.2000 ;
	    RECT 112.6000 107.1000 113.0000 107.2000 ;
	    RECT 92.6000 106.8000 99.3000 107.1000 ;
	    RECT 105.4000 106.8000 113.0000 107.1000 ;
	    RECT 116.6000 107.1000 117.0000 107.2000 ;
	    RECT 122.2000 107.1000 122.6000 107.2000 ;
	    RECT 116.6000 106.8000 122.6000 107.1000 ;
	    RECT 128.6000 107.1000 129.0000 107.2000 ;
	    RECT 131.0000 107.1000 131.4000 107.2000 ;
	    RECT 128.6000 106.8000 131.4000 107.1000 ;
	    RECT 138.2000 106.8000 138.6000 107.2000 ;
	    RECT 41.4000 106.2000 41.7000 106.8000 ;
	    RECT 99.0000 106.2000 99.3000 106.8000 ;
	    RECT 8.6000 106.1000 9.0000 106.2000 ;
	    RECT 14.2000 106.1000 14.6000 106.2000 ;
	    RECT 8.6000 105.8000 14.6000 106.1000 ;
	    RECT 25.4000 105.8000 28.9000 106.1000 ;
	    RECT 41.4000 105.8000 41.8000 106.2000 ;
	    RECT 43.0000 106.1000 43.4000 106.2000 ;
	    RECT 45.4000 106.1000 45.8000 106.2000 ;
	    RECT 43.0000 105.8000 45.8000 106.1000 ;
	    RECT 59.0000 106.1000 59.4000 106.2000 ;
	    RECT 62.2000 106.1000 62.6000 106.2000 ;
	    RECT 65.4000 106.1000 65.8000 106.2000 ;
	    RECT 59.0000 105.8000 65.8000 106.1000 ;
	    RECT 67.0000 105.8000 67.4000 106.2000 ;
	    RECT 79.8000 106.1000 80.2000 106.2000 ;
	    RECT 72.6000 105.8000 80.2000 106.1000 ;
	    RECT 99.0000 105.8000 99.4000 106.2000 ;
	    RECT 113.4000 106.1000 113.8000 106.2000 ;
	    RECT 116.6000 106.1000 117.0000 106.2000 ;
	    RECT 129.4000 106.1000 129.8000 106.2000 ;
	    RECT 135.0000 106.1000 135.4000 106.2000 ;
	    RECT 113.4000 105.8000 135.4000 106.1000 ;
	    RECT 137.4000 106.1000 137.8000 106.2000 ;
	    RECT 141.4000 106.1000 141.8000 106.2000 ;
	    RECT 137.4000 105.8000 141.8000 106.1000 ;
	    RECT 25.4000 105.2000 25.7000 105.8000 ;
	    RECT 28.6000 105.2000 28.9000 105.8000 ;
	    RECT 25.4000 104.8000 25.8000 105.2000 ;
	    RECT 28.6000 104.8000 29.0000 105.2000 ;
	    RECT 43.8000 105.1000 44.2000 105.2000 ;
	    RECT 56.6000 105.1000 57.0000 105.2000 ;
	    RECT 59.0000 105.1000 59.4000 105.2000 ;
	    RECT 43.8000 104.8000 59.4000 105.1000 ;
	    RECT 63.8000 105.1000 64.2000 105.2000 ;
	    RECT 64.6000 105.1000 65.0000 105.2000 ;
	    RECT 63.8000 104.8000 65.0000 105.1000 ;
	    RECT 67.0000 105.1000 67.3000 105.8000 ;
	    RECT 72.6000 105.2000 72.9000 105.8000 ;
	    RECT 67.8000 105.1000 68.2000 105.2000 ;
	    RECT 67.0000 104.8000 68.2000 105.1000 ;
	    RECT 72.6000 104.8000 73.0000 105.2000 ;
	    RECT 96.6000 105.1000 97.0000 105.2000 ;
	    RECT 109.4000 105.1000 109.8000 105.2000 ;
	    RECT 117.4000 105.1000 117.8000 105.2000 ;
	    RECT 96.6000 104.8000 117.8000 105.1000 ;
	    RECT 120.6000 105.1000 121.0000 105.2000 ;
	    RECT 121.4000 105.1000 121.8000 105.2000 ;
	    RECT 127.0000 105.1000 127.4000 105.2000 ;
	    RECT 131.8000 105.1000 132.2000 105.2000 ;
	    RECT 135.8000 105.1000 136.2000 105.2000 ;
	    RECT 120.6000 104.8000 136.2000 105.1000 ;
	    RECT 33.4000 104.1000 33.8000 104.2000 ;
	    RECT 44.6000 104.1000 45.0000 104.2000 ;
	    RECT 33.4000 103.8000 45.0000 104.1000 ;
	    RECT 120.6000 104.1000 121.0000 104.2000 ;
	    RECT 130.2000 104.1000 130.6000 104.2000 ;
	    RECT 146.2000 104.1000 146.6000 104.2000 ;
	    RECT 120.6000 103.8000 128.9000 104.1000 ;
	    RECT 130.2000 103.8000 146.6000 104.1000 ;
	    RECT 128.6000 103.2000 128.9000 103.8000 ;
	    RECT 128.6000 102.8000 129.0000 103.2000 ;
	    RECT 68.6000 100.1000 69.0000 100.2000 ;
	    RECT 81.4000 100.1000 81.8000 100.2000 ;
	    RECT 84.6000 100.1000 85.0000 100.2000 ;
	    RECT 68.6000 99.8000 85.0000 100.1000 ;
	    RECT 125.4000 97.8000 125.8000 98.2000 ;
	    RECT 133.4000 98.1000 133.8000 98.2000 ;
	    RECT 139.8000 98.1000 140.2000 98.2000 ;
	    RECT 133.4000 97.8000 140.2000 98.1000 ;
	    RECT 2.2000 97.1000 2.6000 97.2000 ;
	    RECT 14.2000 97.1000 14.6000 97.2000 ;
	    RECT 19.0000 97.1000 19.4000 97.2000 ;
	    RECT 24.6000 97.1000 25.0000 97.2000 ;
	    RECT 2.2000 96.8000 25.0000 97.1000 ;
	    RECT 39.8000 97.1000 40.2000 97.2000 ;
	    RECT 43.0000 97.1000 43.4000 97.2000 ;
	    RECT 39.8000 96.8000 43.4000 97.1000 ;
	    RECT 59.0000 97.1000 59.4000 97.2000 ;
	    RECT 90.2000 97.1000 90.6000 97.2000 ;
	    RECT 111.0000 97.1000 111.4000 97.2000 ;
	    RECT 59.0000 96.8000 64.9000 97.1000 ;
	    RECT 90.2000 96.8000 111.4000 97.1000 ;
	    RECT 115.8000 97.1000 116.2000 97.2000 ;
	    RECT 119.0000 97.1000 119.4000 97.2000 ;
	    RECT 115.8000 96.8000 119.4000 97.1000 ;
	    RECT 123.8000 97.1000 124.2000 97.2000 ;
	    RECT 125.4000 97.1000 125.7000 97.8000 ;
	    RECT 123.8000 96.8000 125.7000 97.1000 ;
	    RECT 137.4000 97.1000 137.8000 97.2000 ;
	    RECT 140.6000 97.1000 141.0000 97.2000 ;
	    RECT 137.4000 96.8000 141.0000 97.1000 ;
	    RECT 64.6000 96.2000 64.9000 96.8000 ;
	    RECT 21.4000 95.8000 21.8000 96.2000 ;
	    RECT 26.2000 95.8000 26.6000 96.2000 ;
	    RECT 31.8000 96.1000 32.2000 96.2000 ;
	    RECT 43.8000 96.1000 44.2000 96.2000 ;
	    RECT 31.8000 95.8000 44.2000 96.1000 ;
	    RECT 57.4000 96.1000 57.8000 96.2000 ;
	    RECT 63.0000 96.1000 63.4000 96.2000 ;
	    RECT 57.4000 95.8000 63.4000 96.1000 ;
	    RECT 64.6000 95.8000 65.0000 96.2000 ;
	    RECT 75.0000 95.8000 75.4000 96.2000 ;
	    RECT 91.0000 95.8000 91.4000 96.2000 ;
	    RECT 117.4000 96.1000 117.8000 96.2000 ;
	    RECT 119.0000 96.1000 119.4000 96.2000 ;
	    RECT 136.6000 96.1000 137.0000 96.2000 ;
	    RECT 117.4000 95.8000 137.0000 96.1000 ;
	    RECT 13.4000 94.8000 13.8000 95.2000 ;
	    RECT 21.4000 95.1000 21.7000 95.8000 ;
	    RECT 26.2000 95.1000 26.5000 95.8000 ;
	    RECT 21.4000 94.8000 26.5000 95.1000 ;
	    RECT 29.4000 94.8000 29.8000 95.2000 ;
	    RECT 31.8000 95.1000 32.2000 95.2000 ;
	    RECT 32.6000 95.1000 33.0000 95.2000 ;
	    RECT 31.8000 94.8000 33.0000 95.1000 ;
	    RECT 35.8000 95.1000 36.2000 95.2000 ;
	    RECT 45.4000 95.1000 45.8000 95.2000 ;
	    RECT 51.0000 95.1000 51.4000 95.2000 ;
	    RECT 35.8000 94.8000 51.4000 95.1000 ;
	    RECT 55.0000 95.1000 55.4000 95.2000 ;
	    RECT 62.2000 95.1000 62.6000 95.2000 ;
	    RECT 55.0000 94.8000 62.6000 95.1000 ;
	    RECT 63.0000 95.1000 63.4000 95.2000 ;
	    RECT 67.8000 95.1000 68.2000 95.2000 ;
	    RECT 63.0000 94.8000 68.2000 95.1000 ;
	    RECT 71.0000 95.1000 71.4000 95.2000 ;
	    RECT 75.0000 95.1000 75.3000 95.8000 ;
	    RECT 71.0000 94.8000 75.3000 95.1000 ;
	    RECT 91.0000 95.1000 91.3000 95.8000 ;
	    RECT 94.2000 95.1000 94.6000 95.2000 ;
	    RECT 115.0000 95.1000 115.4000 95.2000 ;
	    RECT 91.0000 94.8000 115.4000 95.1000 ;
	    RECT 116.6000 95.1000 117.0000 95.2000 ;
	    RECT 121.4000 95.1000 121.8000 95.2000 ;
	    RECT 116.6000 94.8000 121.8000 95.1000 ;
	    RECT 126.2000 95.1000 126.6000 95.2000 ;
	    RECT 139.8000 95.1000 140.2000 95.2000 ;
	    RECT 126.2000 94.8000 140.2000 95.1000 ;
	    RECT 143.0000 94.8000 143.4000 95.2000 ;
	    RECT 13.4000 94.1000 13.7000 94.8000 ;
	    RECT 18.2000 94.1000 18.6000 94.2000 ;
	    RECT 13.4000 93.8000 18.6000 94.1000 ;
	    RECT 29.4000 94.1000 29.7000 94.8000 ;
	    RECT 32.6000 94.1000 33.0000 94.2000 ;
	    RECT 43.0000 94.1000 43.4000 94.2000 ;
	    RECT 29.4000 93.8000 33.0000 94.1000 ;
	    RECT 35.8000 93.8000 43.4000 94.1000 ;
	    RECT 52.6000 93.8000 53.0000 94.2000 ;
	    RECT 55.8000 93.8000 56.2000 94.2000 ;
	    RECT 67.8000 94.1000 68.2000 94.2000 ;
	    RECT 82.2000 94.1000 82.6000 94.2000 ;
	    RECT 67.8000 93.8000 82.6000 94.1000 ;
	    RECT 85.4000 94.1000 85.8000 94.2000 ;
	    RECT 86.2000 94.1000 86.6000 94.2000 ;
	    RECT 89.4000 94.1000 89.8000 94.2000 ;
	    RECT 91.8000 94.1000 92.2000 94.2000 ;
	    RECT 113.4000 94.1000 113.8000 94.2000 ;
	    RECT 123.8000 94.1000 124.2000 94.2000 ;
	    RECT 85.4000 93.8000 92.2000 94.1000 ;
	    RECT 112.6000 93.8000 124.2000 94.1000 ;
	    RECT 127.0000 94.1000 127.4000 94.2000 ;
	    RECT 138.2000 94.1000 138.6000 94.2000 ;
	    RECT 143.0000 94.1000 143.3000 94.8000 ;
	    RECT 127.0000 93.8000 138.6000 94.1000 ;
	    RECT 139.0000 93.8000 143.3000 94.1000 ;
	    RECT 35.8000 93.2000 36.1000 93.8000 ;
	    RECT 35.8000 92.8000 36.2000 93.2000 ;
	    RECT 40.6000 93.1000 41.0000 93.2000 ;
	    RECT 52.6000 93.1000 52.9000 93.8000 ;
	    RECT 40.6000 92.8000 52.9000 93.1000 ;
	    RECT 55.8000 93.1000 56.1000 93.8000 ;
	    RECT 139.0000 93.2000 139.3000 93.8000 ;
	    RECT 57.4000 93.1000 57.8000 93.2000 ;
	    RECT 55.8000 92.8000 57.8000 93.1000 ;
	    RECT 62.2000 93.1000 62.6000 93.2000 ;
	    RECT 70.2000 93.1000 70.6000 93.2000 ;
	    RECT 62.2000 92.8000 70.6000 93.1000 ;
	    RECT 97.4000 93.1000 97.8000 93.2000 ;
	    RECT 125.4000 93.1000 125.8000 93.2000 ;
	    RECT 97.4000 92.8000 125.8000 93.1000 ;
	    RECT 139.0000 92.8000 139.4000 93.2000 ;
	    RECT 143.0000 93.1000 143.4000 93.2000 ;
	    RECT 144.6000 93.1000 145.0000 93.2000 ;
	    RECT 143.0000 92.8000 145.0000 93.1000 ;
	    RECT 11.8000 92.1000 12.2000 92.2000 ;
	    RECT 14.2000 92.1000 14.6000 92.2000 ;
	    RECT 11.8000 91.8000 14.6000 92.1000 ;
	    RECT 27.0000 92.1000 27.4000 92.2000 ;
	    RECT 30.2000 92.1000 30.6000 92.2000 ;
	    RECT 27.0000 91.8000 30.6000 92.1000 ;
	    RECT 41.4000 92.1000 41.8000 92.2000 ;
	    RECT 53.4000 92.1000 53.8000 92.2000 ;
	    RECT 58.2000 92.1000 58.6000 92.2000 ;
	    RECT 41.4000 91.8000 58.6000 92.1000 ;
	    RECT 96.6000 92.1000 97.0000 92.2000 ;
	    RECT 117.4000 92.1000 117.8000 92.2000 ;
	    RECT 124.6000 92.1000 125.0000 92.2000 ;
	    RECT 130.2000 92.1000 130.6000 92.2000 ;
	    RECT 96.6000 91.8000 117.8000 92.1000 ;
	    RECT 123.8000 91.8000 130.6000 92.1000 ;
	    RECT 24.6000 91.1000 25.0000 91.2000 ;
	    RECT 33.4000 91.1000 33.8000 91.2000 ;
	    RECT 24.6000 90.8000 33.8000 91.1000 ;
	    RECT 103.0000 91.1000 103.4000 91.2000 ;
	    RECT 105.4000 91.1000 105.8000 91.2000 ;
	    RECT 103.0000 90.8000 105.8000 91.1000 ;
	    RECT 115.0000 91.1000 115.4000 91.2000 ;
	    RECT 116.6000 91.1000 117.0000 91.2000 ;
	    RECT 115.0000 90.8000 117.0000 91.1000 ;
	    RECT 15.0000 90.1000 15.4000 90.2000 ;
	    RECT 15.8000 90.1000 16.2000 90.2000 ;
	    RECT 71.8000 90.1000 72.2000 90.2000 ;
	    RECT 72.6000 90.1000 73.0000 90.2000 ;
	    RECT 15.0000 89.8000 73.0000 90.1000 ;
	    RECT 112.6000 90.1000 113.0000 90.2000 ;
	    RECT 114.2000 90.1000 114.6000 90.2000 ;
	    RECT 121.4000 90.1000 121.8000 90.2000 ;
	    RECT 112.6000 89.8000 121.8000 90.1000 ;
	    RECT 4.6000 89.1000 5.0000 89.2000 ;
	    RECT 28.6000 89.1000 29.0000 89.2000 ;
	    RECT 46.2000 89.1000 46.6000 89.2000 ;
	    RECT 53.4000 89.1000 53.8000 89.2000 ;
	    RECT 56.6000 89.1000 57.0000 89.2000 ;
	    RECT 62.2000 89.1000 62.6000 89.2000 ;
	    RECT 4.6000 88.8000 57.0000 89.1000 ;
	    RECT 57.4000 88.8000 62.6000 89.1000 ;
	    RECT 75.0000 89.1000 75.4000 89.2000 ;
	    RECT 83.8000 89.1000 84.2000 89.2000 ;
	    RECT 75.0000 88.8000 84.2000 89.1000 ;
	    RECT 87.0000 89.1000 87.4000 89.2000 ;
	    RECT 87.8000 89.1000 88.2000 89.2000 ;
	    RECT 87.0000 88.8000 88.2000 89.1000 ;
	    RECT 108.6000 89.1000 109.0000 89.2000 ;
	    RECT 115.0000 89.1000 115.4000 89.2000 ;
	    RECT 108.6000 88.8000 115.4000 89.1000 ;
	    RECT 12.6000 87.8000 13.0000 88.2000 ;
	    RECT 35.0000 87.8000 35.4000 88.2000 ;
	    RECT 51.0000 88.1000 51.4000 88.2000 ;
	    RECT 57.4000 88.1000 57.7000 88.8000 ;
	    RECT 51.0000 87.8000 57.7000 88.1000 ;
	    RECT 59.8000 88.1000 60.2000 88.2000 ;
	    RECT 64.6000 88.1000 65.0000 88.2000 ;
	    RECT 77.4000 88.1000 77.8000 88.2000 ;
	    RECT 59.8000 87.8000 77.8000 88.1000 ;
	    RECT 78.2000 88.1000 78.6000 88.2000 ;
	    RECT 86.2000 88.1000 86.6000 88.2000 ;
	    RECT 78.2000 87.8000 86.6000 88.1000 ;
	    RECT 93.4000 88.1000 93.8000 88.2000 ;
	    RECT 95.0000 88.1000 95.4000 88.2000 ;
	    RECT 93.4000 87.8000 95.4000 88.1000 ;
	    RECT 6.2000 87.1000 6.6000 87.2000 ;
	    RECT 12.6000 87.1000 12.9000 87.8000 ;
	    RECT 6.2000 86.8000 12.9000 87.1000 ;
	    RECT 17.4000 87.1000 17.8000 87.2000 ;
	    RECT 23.0000 87.1000 23.4000 87.2000 ;
	    RECT 35.0000 87.1000 35.3000 87.8000 ;
	    RECT 47.0000 87.1000 47.4000 87.2000 ;
	    RECT 17.4000 86.8000 18.5000 87.1000 ;
	    RECT 23.0000 86.8000 35.3000 87.1000 ;
	    RECT 35.8000 86.8000 47.4000 87.1000 ;
	    RECT 57.4000 86.8000 57.8000 87.2000 ;
	    RECT 64.6000 87.1000 65.0000 87.2000 ;
	    RECT 65.4000 87.1000 65.8000 87.2000 ;
	    RECT 64.6000 86.8000 65.8000 87.1000 ;
	    RECT 69.4000 87.1000 69.8000 87.2000 ;
	    RECT 71.8000 87.1000 72.2000 87.2000 ;
	    RECT 69.4000 86.8000 72.2000 87.1000 ;
	    RECT 86.2000 87.1000 86.5000 87.8000 ;
	    RECT 95.0000 87.1000 95.4000 87.2000 ;
	    RECT 86.2000 86.8000 95.4000 87.1000 ;
	    RECT 107.0000 87.1000 107.4000 87.2000 ;
	    RECT 109.4000 87.1000 109.8000 87.2000 ;
	    RECT 107.0000 86.8000 109.8000 87.1000 ;
	    RECT 119.0000 87.1000 119.4000 87.2000 ;
	    RECT 119.8000 87.1000 120.2000 87.2000 ;
	    RECT 119.0000 86.8000 120.2000 87.1000 ;
	    RECT 18.2000 86.2000 18.5000 86.8000 ;
	    RECT 18.2000 86.1000 18.6000 86.2000 ;
	    RECT 24.6000 86.1000 25.0000 86.2000 ;
	    RECT 18.2000 85.8000 25.0000 86.1000 ;
	    RECT 33.4000 86.1000 33.8000 86.2000 ;
	    RECT 35.8000 86.1000 36.1000 86.8000 ;
	    RECT 33.4000 85.8000 36.1000 86.1000 ;
	    RECT 43.0000 86.1000 43.4000 86.2000 ;
	    RECT 44.6000 86.1000 45.0000 86.2000 ;
	    RECT 43.0000 85.8000 45.0000 86.1000 ;
	    RECT 48.6000 86.1000 49.0000 86.2000 ;
	    RECT 54.2000 86.1000 54.6000 86.2000 ;
	    RECT 48.6000 85.8000 54.6000 86.1000 ;
	    RECT 57.4000 86.1000 57.7000 86.8000 ;
	    RECT 58.2000 86.1000 58.6000 86.2000 ;
	    RECT 57.4000 85.8000 58.6000 86.1000 ;
	    RECT 60.6000 86.1000 61.0000 86.2000 ;
	    RECT 63.0000 86.1000 63.4000 86.2000 ;
	    RECT 60.6000 85.8000 63.4000 86.1000 ;
	    RECT 74.2000 86.1000 74.6000 86.2000 ;
	    RECT 87.8000 86.1000 88.2000 86.2000 ;
	    RECT 108.6000 86.1000 109.0000 86.2000 ;
	    RECT 110.2000 86.1000 110.6000 86.2000 ;
	    RECT 119.0000 86.1000 119.4000 86.2000 ;
	    RECT 131.0000 86.1000 131.4000 86.2000 ;
	    RECT 74.2000 85.8000 88.2000 86.1000 ;
	    RECT 107.8000 85.8000 131.4000 86.1000 ;
	    RECT 21.4000 85.1000 21.8000 85.2000 ;
	    RECT 27.8000 85.1000 28.2000 85.2000 ;
	    RECT 21.4000 84.8000 28.2000 85.1000 ;
	    RECT 45.4000 85.1000 45.8000 85.2000 ;
	    RECT 49.4000 85.1000 49.8000 85.2000 ;
	    RECT 45.4000 84.8000 49.8000 85.1000 ;
	    RECT 56.6000 85.1000 57.0000 85.2000 ;
	    RECT 58.2000 85.1000 58.6000 85.2000 ;
	    RECT 56.6000 84.8000 58.6000 85.1000 ;
	    RECT 59.0000 85.1000 59.4000 85.2000 ;
	    RECT 65.4000 85.1000 65.8000 85.2000 ;
	    RECT 59.0000 84.8000 65.8000 85.1000 ;
	    RECT 82.2000 85.1000 82.6000 85.2000 ;
	    RECT 95.8000 85.1000 96.2000 85.2000 ;
	    RECT 98.2000 85.1000 98.6000 85.2000 ;
	    RECT 82.2000 84.8000 98.6000 85.1000 ;
	    RECT 110.2000 85.1000 110.6000 85.2000 ;
	    RECT 116.6000 85.1000 117.0000 85.2000 ;
	    RECT 110.2000 84.8000 117.0000 85.1000 ;
	    RECT 9.4000 84.1000 9.8000 84.2000 ;
	    RECT 31.0000 84.1000 31.4000 84.2000 ;
	    RECT 9.4000 83.8000 31.4000 84.1000 ;
	    RECT 34.2000 84.1000 34.6000 84.2000 ;
	    RECT 43.8000 84.1000 44.2000 84.2000 ;
	    RECT 34.2000 83.8000 44.2000 84.1000 ;
	    RECT 53.4000 84.1000 53.8000 84.2000 ;
	    RECT 68.6000 84.1000 69.0000 84.2000 ;
	    RECT 53.4000 83.8000 69.0000 84.1000 ;
	    RECT 93.4000 84.1000 93.8000 84.2000 ;
	    RECT 107.0000 84.1000 107.4000 84.2000 ;
	    RECT 93.4000 83.8000 107.4000 84.1000 ;
	    RECT 108.6000 84.1000 109.0000 84.2000 ;
	    RECT 114.2000 84.1000 114.6000 84.2000 ;
	    RECT 108.6000 83.8000 114.6000 84.1000 ;
	    RECT 119.8000 84.1000 120.2000 84.2000 ;
	    RECT 120.6000 84.1000 121.0000 84.2000 ;
	    RECT 132.6000 84.1000 133.0000 84.2000 ;
	    RECT 142.2000 84.1000 142.6000 84.2000 ;
	    RECT 145.4000 84.1000 145.8000 84.2000 ;
	    RECT 119.8000 83.8000 145.8000 84.1000 ;
	    RECT 13.4000 83.1000 13.8000 83.2000 ;
	    RECT 19.0000 83.1000 19.4000 83.2000 ;
	    RECT 13.4000 82.8000 19.4000 83.1000 ;
	    RECT 43.8000 83.1000 44.2000 83.2000 ;
	    RECT 47.8000 83.1000 48.2000 83.2000 ;
	    RECT 51.8000 83.1000 52.2000 83.2000 ;
	    RECT 43.8000 82.8000 52.2000 83.1000 ;
	    RECT 87.0000 83.1000 87.4000 83.2000 ;
	    RECT 99.0000 83.1000 99.4000 83.2000 ;
	    RECT 87.0000 82.8000 99.4000 83.1000 ;
	    RECT 99.8000 83.1000 100.2000 83.2000 ;
	    RECT 118.2000 83.1000 118.6000 83.2000 ;
	    RECT 99.8000 82.8000 118.6000 83.1000 ;
	    RECT 106.2000 82.1000 106.6000 82.2000 ;
	    RECT 122.2000 82.1000 122.6000 82.2000 ;
	    RECT 106.2000 81.8000 122.6000 82.1000 ;
	    RECT 71.0000 81.1000 71.4000 81.2000 ;
	    RECT 71.8000 81.1000 72.2000 81.2000 ;
	    RECT 71.0000 80.8000 72.2000 81.1000 ;
	    RECT 72.6000 81.1000 73.0000 81.2000 ;
	    RECT 87.8000 81.1000 88.2000 81.2000 ;
	    RECT 143.8000 81.1000 144.2000 81.2000 ;
	    RECT 144.6000 81.1000 145.0000 81.2000 ;
	    RECT 72.6000 80.8000 145.0000 81.1000 ;
	    RECT 109.4000 80.1000 109.8000 80.2000 ;
	    RECT 112.6000 80.1000 113.0000 80.2000 ;
	    RECT 109.4000 79.8000 113.0000 80.1000 ;
	    RECT 129.4000 80.1000 129.8000 80.2000 ;
	    RECT 135.0000 80.1000 135.4000 80.2000 ;
	    RECT 129.4000 79.8000 135.4000 80.1000 ;
	    RECT 62.2000 79.1000 62.6000 79.2000 ;
	    RECT 70.2000 79.1000 70.6000 79.2000 ;
	    RECT 83.0000 79.1000 83.4000 79.2000 ;
	    RECT 62.2000 78.8000 83.4000 79.1000 ;
	    RECT 99.0000 79.1000 99.4000 79.2000 ;
	    RECT 110.2000 79.1000 110.6000 79.2000 ;
	    RECT 99.0000 78.8000 110.6000 79.1000 ;
	    RECT 35.8000 78.1000 36.2000 78.2000 ;
	    RECT 51.0000 78.1000 51.4000 78.2000 ;
	    RECT 35.8000 77.8000 51.4000 78.1000 ;
	    RECT 57.4000 78.1000 57.8000 78.2000 ;
	    RECT 67.8000 78.1000 68.2000 78.2000 ;
	    RECT 57.4000 77.8000 68.2000 78.1000 ;
	    RECT 77.4000 78.1000 77.8000 78.2000 ;
	    RECT 79.0000 78.1000 79.4000 78.2000 ;
	    RECT 83.0000 78.1000 83.4000 78.2000 ;
	    RECT 103.8000 78.1000 104.2000 78.2000 ;
	    RECT 77.4000 77.8000 104.2000 78.1000 ;
	    RECT 108.6000 78.1000 109.0000 78.2000 ;
	    RECT 112.6000 78.1000 113.0000 78.2000 ;
	    RECT 108.6000 77.8000 113.0000 78.1000 ;
	    RECT 114.2000 77.8000 114.6000 78.2000 ;
	    RECT 115.0000 78.1000 115.4000 78.2000 ;
	    RECT 119.8000 78.1000 120.2000 78.2000 ;
	    RECT 115.0000 77.8000 120.2000 78.1000 ;
	    RECT 138.2000 77.8000 138.6000 78.2000 ;
	    RECT 12.6000 77.1000 13.0000 77.2000 ;
	    RECT 24.6000 77.1000 25.0000 77.2000 ;
	    RECT 12.6000 76.8000 25.0000 77.1000 ;
	    RECT 39.0000 76.8000 39.4000 77.2000 ;
	    RECT 40.6000 77.1000 41.0000 77.2000 ;
	    RECT 59.8000 77.1000 60.2000 77.2000 ;
	    RECT 40.6000 76.8000 60.2000 77.1000 ;
	    RECT 81.4000 76.8000 81.8000 77.2000 ;
	    RECT 89.4000 77.1000 89.8000 77.2000 ;
	    RECT 97.4000 77.1000 97.8000 77.2000 ;
	    RECT 89.4000 76.8000 97.8000 77.1000 ;
	    RECT 98.2000 77.1000 98.6000 77.2000 ;
	    RECT 99.0000 77.1000 99.4000 77.2000 ;
	    RECT 107.0000 77.1000 107.4000 77.2000 ;
	    RECT 98.2000 76.8000 107.4000 77.1000 ;
	    RECT 114.2000 77.1000 114.5000 77.8000 ;
	    RECT 122.2000 77.1000 122.6000 77.2000 ;
	    RECT 114.2000 76.8000 122.6000 77.1000 ;
	    RECT 124.6000 77.1000 125.0000 77.2000 ;
	    RECT 130.2000 77.1000 130.6000 77.2000 ;
	    RECT 124.6000 76.8000 130.6000 77.1000 ;
	    RECT 131.8000 77.1000 132.2000 77.2000 ;
	    RECT 138.2000 77.1000 138.5000 77.8000 ;
	    RECT 131.8000 76.8000 138.5000 77.1000 ;
	    RECT 143.0000 77.1000 143.4000 77.2000 ;
	    RECT 145.4000 77.1000 145.8000 77.2000 ;
	    RECT 143.0000 76.8000 145.8000 77.1000 ;
	    RECT 15.8000 76.1000 16.2000 76.2000 ;
	    RECT 16.6000 76.1000 17.0000 76.2000 ;
	    RECT 25.4000 76.1000 25.8000 76.2000 ;
	    RECT 15.8000 75.8000 25.8000 76.1000 ;
	    RECT 31.0000 75.8000 31.4000 76.2000 ;
	    RECT 39.0000 76.1000 39.3000 76.8000 ;
	    RECT 46.2000 76.1000 46.6000 76.2000 ;
	    RECT 39.0000 75.8000 46.6000 76.1000 ;
	    RECT 69.4000 76.1000 69.8000 76.2000 ;
	    RECT 79.8000 76.1000 80.2000 76.2000 ;
	    RECT 69.4000 75.8000 80.2000 76.1000 ;
	    RECT 81.4000 76.1000 81.7000 76.8000 ;
	    RECT 85.4000 76.1000 85.8000 76.2000 ;
	    RECT 88.6000 76.1000 89.0000 76.2000 ;
	    RECT 81.4000 75.8000 89.0000 76.1000 ;
	    RECT 91.0000 76.1000 91.4000 76.2000 ;
	    RECT 103.8000 76.1000 104.2000 76.2000 ;
	    RECT 91.0000 75.8000 104.2000 76.1000 ;
	    RECT 111.8000 76.1000 112.2000 76.2000 ;
	    RECT 115.8000 76.1000 116.2000 76.2000 ;
	    RECT 111.8000 75.8000 116.2000 76.1000 ;
	    RECT 116.6000 76.1000 117.0000 76.2000 ;
	    RECT 125.4000 76.1000 125.8000 76.2000 ;
	    RECT 137.4000 76.1000 137.8000 76.2000 ;
	    RECT 116.6000 75.8000 125.8000 76.1000 ;
	    RECT 136.6000 75.8000 137.8000 76.1000 ;
	    RECT 7.0000 75.1000 7.4000 75.2000 ;
	    RECT 13.4000 75.1000 13.8000 75.2000 ;
	    RECT 30.2000 75.1000 30.6000 75.2000 ;
	    RECT 7.0000 74.8000 13.8000 75.1000 ;
	    RECT 29.4000 74.8000 30.6000 75.1000 ;
	    RECT 31.0000 75.1000 31.3000 75.8000 ;
	    RECT 136.6000 75.2000 136.9000 75.8000 ;
	    RECT 42.2000 75.1000 42.6000 75.2000 ;
	    RECT 31.0000 74.8000 42.6000 75.1000 ;
	    RECT 51.8000 75.1000 52.2000 75.2000 ;
	    RECT 56.6000 75.1000 57.0000 75.2000 ;
	    RECT 66.2000 75.1000 66.6000 75.2000 ;
	    RECT 51.8000 74.8000 66.6000 75.1000 ;
	    RECT 84.6000 75.1000 85.0000 75.2000 ;
	    RECT 88.6000 75.1000 89.0000 75.2000 ;
	    RECT 84.6000 74.8000 89.0000 75.1000 ;
	    RECT 91.0000 75.1000 91.4000 75.2000 ;
	    RECT 113.4000 75.1000 113.8000 75.2000 ;
	    RECT 115.8000 75.1000 116.2000 75.2000 ;
	    RECT 116.6000 75.1000 117.0000 75.2000 ;
	    RECT 91.0000 74.8000 117.0000 75.1000 ;
	    RECT 123.0000 75.1000 123.4000 75.2000 ;
	    RECT 126.2000 75.1000 126.6000 75.2000 ;
	    RECT 123.0000 74.8000 126.6000 75.1000 ;
	    RECT 136.6000 74.8000 137.0000 75.2000 ;
	    RECT 138.2000 75.1000 138.6000 75.2000 ;
	    RECT 139.8000 75.1000 140.2000 75.2000 ;
	    RECT 142.2000 75.1000 142.6000 75.2000 ;
	    RECT 138.2000 74.8000 142.6000 75.1000 ;
	    RECT 6.2000 74.1000 6.6000 74.2000 ;
	    RECT 11.8000 74.1000 12.2000 74.2000 ;
	    RECT 18.2000 74.1000 18.6000 74.2000 ;
	    RECT 6.2000 73.8000 18.6000 74.1000 ;
	    RECT 23.8000 74.1000 24.2000 74.2000 ;
	    RECT 27.8000 74.1000 28.2000 74.2000 ;
	    RECT 23.8000 73.8000 28.2000 74.1000 ;
	    RECT 37.4000 74.1000 37.8000 74.2000 ;
	    RECT 39.8000 74.1000 40.2000 74.2000 ;
	    RECT 37.4000 73.8000 40.2000 74.1000 ;
	    RECT 43.0000 74.1000 43.4000 74.2000 ;
	    RECT 46.2000 74.1000 46.6000 74.2000 ;
	    RECT 43.0000 73.8000 46.6000 74.1000 ;
	    RECT 50.2000 74.1000 50.6000 74.2000 ;
	    RECT 55.0000 74.1000 55.4000 74.2000 ;
	    RECT 50.2000 73.8000 55.4000 74.1000 ;
	    RECT 89.4000 74.1000 89.8000 74.2000 ;
	    RECT 91.8000 74.1000 92.2000 74.2000 ;
	    RECT 89.4000 73.8000 92.2000 74.1000 ;
	    RECT 103.8000 74.1000 104.2000 74.2000 ;
	    RECT 119.0000 74.1000 119.4000 74.2000 ;
	    RECT 143.8000 74.1000 144.2000 74.2000 ;
	    RECT 103.8000 73.8000 144.2000 74.1000 ;
	    RECT 3.8000 73.1000 4.2000 73.2000 ;
	    RECT 5.4000 73.1000 5.8000 73.2000 ;
	    RECT 3.8000 72.8000 5.8000 73.1000 ;
	    RECT 9.4000 73.1000 9.8000 73.2000 ;
	    RECT 15.8000 73.1000 16.2000 73.2000 ;
	    RECT 9.4000 72.8000 16.2000 73.1000 ;
	    RECT 20.6000 73.1000 21.0000 73.2000 ;
	    RECT 23.0000 73.1000 23.4000 73.2000 ;
	    RECT 20.6000 72.8000 23.4000 73.1000 ;
	    RECT 24.6000 73.1000 25.0000 73.2000 ;
	    RECT 25.4000 73.1000 25.8000 73.2000 ;
	    RECT 24.6000 72.8000 25.8000 73.1000 ;
	    RECT 27.8000 73.1000 28.1000 73.8000 ;
	    RECT 28.6000 73.1000 29.0000 73.2000 ;
	    RECT 29.4000 73.1000 29.8000 73.2000 ;
	    RECT 31.0000 73.1000 31.4000 73.2000 ;
	    RECT 27.8000 72.8000 31.4000 73.1000 ;
	    RECT 36.6000 73.1000 37.0000 73.2000 ;
	    RECT 39.8000 73.1000 40.2000 73.2000 ;
	    RECT 36.6000 72.8000 40.2000 73.1000 ;
	    RECT 45.4000 73.1000 45.8000 73.2000 ;
	    RECT 54.2000 73.1000 54.6000 73.2000 ;
	    RECT 45.4000 72.8000 54.6000 73.1000 ;
	    RECT 79.0000 73.1000 79.4000 73.2000 ;
	    RECT 81.4000 73.1000 81.8000 73.2000 ;
	    RECT 79.0000 72.8000 81.8000 73.1000 ;
	    RECT 96.6000 73.1000 97.0000 73.2000 ;
	    RECT 108.6000 73.1000 109.0000 73.2000 ;
	    RECT 114.2000 73.1000 114.6000 73.2000 ;
	    RECT 96.6000 72.8000 114.6000 73.1000 ;
	    RECT 115.8000 73.1000 116.2000 73.2000 ;
	    RECT 118.2000 73.1000 118.6000 73.2000 ;
	    RECT 115.8000 72.8000 118.6000 73.1000 ;
	    RECT 123.0000 73.1000 123.4000 73.2000 ;
	    RECT 126.2000 73.1000 126.6000 73.2000 ;
	    RECT 123.0000 72.8000 126.6000 73.1000 ;
	    RECT 130.2000 73.1000 130.6000 73.2000 ;
	    RECT 137.4000 73.1000 137.8000 73.2000 ;
	    RECT 139.8000 73.1000 140.2000 73.2000 ;
	    RECT 130.2000 72.8000 140.2000 73.1000 ;
	    RECT 10.2000 72.1000 10.6000 72.2000 ;
	    RECT 12.6000 72.1000 13.0000 72.2000 ;
	    RECT 10.2000 71.8000 13.0000 72.1000 ;
	    RECT 25.4000 72.1000 25.8000 72.2000 ;
	    RECT 31.8000 72.1000 32.2000 72.2000 ;
	    RECT 32.6000 72.1000 33.0000 72.2000 ;
	    RECT 38.2000 72.1000 38.6000 72.2000 ;
	    RECT 25.4000 71.8000 38.6000 72.1000 ;
	    RECT 48.6000 72.1000 49.0000 72.2000 ;
	    RECT 51.8000 72.1000 52.2000 72.2000 ;
	    RECT 48.6000 71.8000 52.2000 72.1000 ;
	    RECT 71.0000 72.1000 71.4000 72.2000 ;
	    RECT 72.6000 72.1000 73.0000 72.2000 ;
	    RECT 71.0000 71.8000 73.0000 72.1000 ;
	    RECT 81.4000 72.1000 81.8000 72.2000 ;
	    RECT 94.2000 72.1000 94.6000 72.2000 ;
	    RECT 96.6000 72.1000 97.0000 72.2000 ;
	    RECT 81.4000 71.8000 97.0000 72.1000 ;
	    RECT 97.4000 72.1000 97.8000 72.2000 ;
	    RECT 113.4000 72.1000 113.8000 72.2000 ;
	    RECT 97.4000 71.8000 113.8000 72.1000 ;
	    RECT 127.0000 72.1000 127.4000 72.2000 ;
	    RECT 134.2000 72.1000 134.6000 72.2000 ;
	    RECT 127.0000 71.8000 134.6000 72.1000 ;
	    RECT 135.0000 72.1000 135.4000 72.2000 ;
	    RECT 137.4000 72.1000 137.8000 72.2000 ;
	    RECT 135.0000 71.8000 137.8000 72.1000 ;
	    RECT 72.6000 71.1000 73.0000 71.2000 ;
	    RECT 91.0000 71.1000 91.4000 71.2000 ;
	    RECT 72.6000 70.8000 91.4000 71.1000 ;
	    RECT 105.4000 71.1000 105.8000 71.2000 ;
	    RECT 116.6000 71.1000 117.0000 71.2000 ;
	    RECT 105.4000 70.8000 117.0000 71.1000 ;
	    RECT 117.4000 71.1000 117.8000 71.2000 ;
	    RECT 127.8000 71.1000 128.2000 71.2000 ;
	    RECT 117.4000 70.8000 128.2000 71.1000 ;
	    RECT 133.4000 71.1000 133.8000 71.2000 ;
	    RECT 136.6000 71.1000 137.0000 71.2000 ;
	    RECT 133.4000 70.8000 137.0000 71.1000 ;
	    RECT 17.4000 70.1000 17.8000 70.2000 ;
	    RECT 20.6000 70.1000 21.0000 70.2000 ;
	    RECT 17.4000 69.8000 21.0000 70.1000 ;
	    RECT 54.2000 70.1000 54.6000 70.2000 ;
	    RECT 59.0000 70.1000 59.4000 70.2000 ;
	    RECT 54.2000 69.8000 59.4000 70.1000 ;
	    RECT 76.6000 70.1000 77.0000 70.2000 ;
	    RECT 80.6000 70.1000 81.0000 70.2000 ;
	    RECT 83.0000 70.1000 83.4000 70.2000 ;
	    RECT 84.6000 70.1000 85.0000 70.2000 ;
	    RECT 76.6000 69.8000 85.0000 70.1000 ;
	    RECT 86.2000 70.1000 86.6000 70.2000 ;
	    RECT 109.4000 70.1000 109.8000 70.2000 ;
	    RECT 112.6000 70.1000 113.0000 70.2000 ;
	    RECT 133.4000 70.1000 133.8000 70.2000 ;
	    RECT 86.2000 69.8000 95.3000 70.1000 ;
	    RECT 109.4000 69.8000 133.8000 70.1000 ;
	    RECT 7.0000 69.1000 7.4000 69.2000 ;
	    RECT 25.4000 69.1000 25.8000 69.2000 ;
	    RECT 27.0000 69.1000 27.4000 69.2000 ;
	    RECT 7.0000 68.8000 27.4000 69.1000 ;
	    RECT 55.0000 69.1000 55.4000 69.2000 ;
	    RECT 60.6000 69.1000 61.0000 69.2000 ;
	    RECT 55.0000 68.8000 61.0000 69.1000 ;
	    RECT 87.0000 69.1000 87.4000 69.2000 ;
	    RECT 90.2000 69.1000 90.6000 69.2000 ;
	    RECT 87.0000 68.8000 90.6000 69.1000 ;
	    RECT 91.0000 69.1000 91.4000 69.2000 ;
	    RECT 94.2000 69.1000 94.6000 69.2000 ;
	    RECT 91.0000 68.8000 94.6000 69.1000 ;
	    RECT 95.0000 69.1000 95.3000 69.8000 ;
	    RECT 100.6000 69.1000 101.0000 69.2000 ;
	    RECT 95.0000 68.8000 101.0000 69.1000 ;
	    RECT 124.6000 68.8000 125.0000 69.2000 ;
	    RECT 135.8000 69.1000 136.2000 69.2000 ;
	    RECT 135.8000 68.8000 139.3000 69.1000 ;
	    RECT 12.6000 67.8000 13.0000 68.2000 ;
	    RECT 19.0000 68.1000 19.4000 68.2000 ;
	    RECT 22.2000 68.1000 22.6000 68.2000 ;
	    RECT 19.0000 67.8000 22.6000 68.1000 ;
	    RECT 43.0000 68.1000 43.4000 68.2000 ;
	    RECT 54.2000 68.1000 54.6000 68.2000 ;
	    RECT 70.2000 68.1000 70.6000 68.2000 ;
	    RECT 43.0000 67.8000 70.6000 68.1000 ;
	    RECT 83.8000 68.1000 84.2000 68.2000 ;
	    RECT 86.2000 68.1000 86.6000 68.2000 ;
	    RECT 105.4000 68.1000 105.8000 68.2000 ;
	    RECT 83.8000 67.8000 105.8000 68.1000 ;
	    RECT 124.6000 68.1000 124.9000 68.8000 ;
	    RECT 139.0000 68.2000 139.3000 68.8000 ;
	    RECT 127.8000 68.1000 128.2000 68.2000 ;
	    RECT 124.6000 67.8000 128.2000 68.1000 ;
	    RECT 133.4000 68.1000 133.8000 68.2000 ;
	    RECT 138.2000 68.1000 138.6000 68.2000 ;
	    RECT 133.4000 67.8000 138.6000 68.1000 ;
	    RECT 139.0000 67.8000 139.4000 68.2000 ;
	    RECT 139.8000 67.8000 140.2000 68.2000 ;
	    RECT 3.8000 67.1000 4.2000 67.2000 ;
	    RECT 12.6000 67.1000 12.9000 67.8000 ;
	    RECT 3.8000 66.8000 12.9000 67.1000 ;
	    RECT 14.2000 67.1000 14.6000 67.2000 ;
	    RECT 27.8000 67.1000 28.2000 67.2000 ;
	    RECT 32.6000 67.1000 33.0000 67.2000 ;
	    RECT 14.2000 66.8000 33.0000 67.1000 ;
	    RECT 33.4000 67.1000 33.8000 67.2000 ;
	    RECT 37.4000 67.1000 37.8000 67.2000 ;
	    RECT 33.4000 66.8000 37.8000 67.1000 ;
	    RECT 39.8000 67.1000 40.2000 67.2000 ;
	    RECT 41.4000 67.1000 41.8000 67.2000 ;
	    RECT 43.0000 67.1000 43.4000 67.2000 ;
	    RECT 39.8000 66.8000 43.4000 67.1000 ;
	    RECT 62.2000 67.1000 62.6000 67.2000 ;
	    RECT 64.6000 67.1000 65.0000 67.2000 ;
	    RECT 62.2000 66.8000 65.0000 67.1000 ;
	    RECT 70.2000 66.8000 70.5000 67.8000 ;
	    RECT 79.0000 67.1000 79.4000 67.2000 ;
	    RECT 82.2000 67.1000 82.6000 67.2000 ;
	    RECT 84.6000 67.1000 85.0000 67.2000 ;
	    RECT 89.4000 67.1000 89.8000 67.2000 ;
	    RECT 79.0000 66.8000 89.8000 67.1000 ;
	    RECT 90.2000 67.1000 90.6000 67.2000 ;
	    RECT 92.6000 67.1000 93.0000 67.2000 ;
	    RECT 90.2000 66.8000 93.0000 67.1000 ;
	    RECT 95.8000 66.8000 96.2000 67.2000 ;
	    RECT 111.8000 67.1000 112.2000 67.2000 ;
	    RECT 123.0000 67.1000 123.4000 67.2000 ;
	    RECT 111.8000 66.8000 123.4000 67.1000 ;
	    RECT 124.6000 67.1000 125.0000 67.2000 ;
	    RECT 125.4000 67.1000 125.8000 67.2000 ;
	    RECT 130.2000 67.1000 130.6000 67.2000 ;
	    RECT 124.6000 66.8000 130.6000 67.1000 ;
	    RECT 132.6000 67.1000 133.0000 67.2000 ;
	    RECT 139.8000 67.1000 140.1000 67.8000 ;
	    RECT 132.6000 66.8000 140.1000 67.1000 ;
	    RECT 20.6000 66.1000 21.0000 66.2000 ;
	    RECT 25.4000 66.1000 25.8000 66.2000 ;
	    RECT 35.8000 66.1000 36.2000 66.2000 ;
	    RECT 9.4000 65.8000 16.1000 66.1000 ;
	    RECT 20.6000 65.8000 36.2000 66.1000 ;
	    RECT 40.6000 66.1000 41.0000 66.2000 ;
	    RECT 55.0000 66.1000 55.4000 66.2000 ;
	    RECT 40.6000 65.8000 55.4000 66.1000 ;
	    RECT 70.2000 66.1000 70.6000 66.2000 ;
	    RECT 71.0000 66.1000 71.4000 66.2000 ;
	    RECT 70.2000 65.8000 71.4000 66.1000 ;
	    RECT 81.4000 66.1000 81.8000 66.2000 ;
	    RECT 85.4000 66.1000 85.8000 66.2000 ;
	    RECT 90.2000 66.1000 90.6000 66.2000 ;
	    RECT 81.4000 65.8000 90.6000 66.1000 ;
	    RECT 95.8000 66.1000 96.1000 66.8000 ;
	    RECT 105.4000 66.1000 105.8000 66.2000 ;
	    RECT 95.8000 65.8000 105.8000 66.1000 ;
	    RECT 109.4000 65.8000 109.8000 66.2000 ;
	    RECT 112.6000 66.1000 113.0000 66.2000 ;
	    RECT 115.8000 66.1000 116.2000 66.2000 ;
	    RECT 112.6000 65.8000 116.2000 66.1000 ;
	    RECT 117.4000 65.8000 117.8000 66.2000 ;
	    RECT 120.6000 66.1000 121.0000 66.2000 ;
	    RECT 125.4000 66.1000 125.8000 66.2000 ;
	    RECT 127.0000 66.1000 127.4000 66.2000 ;
	    RECT 128.6000 66.1000 129.0000 66.2000 ;
	    RECT 120.6000 65.8000 127.4000 66.1000 ;
	    RECT 127.8000 65.8000 129.0000 66.1000 ;
	    RECT 133.4000 66.1000 133.8000 66.2000 ;
	    RECT 135.8000 66.1000 136.2000 66.2000 ;
	    RECT 133.4000 65.8000 136.2000 66.1000 ;
	    RECT 138.2000 66.1000 138.6000 66.2000 ;
	    RECT 140.6000 66.1000 141.0000 66.2000 ;
	    RECT 138.2000 65.8000 141.0000 66.1000 ;
	    RECT 9.4000 65.2000 9.7000 65.8000 ;
	    RECT 15.8000 65.2000 16.1000 65.8000 ;
	    RECT 9.4000 64.8000 9.8000 65.2000 ;
	    RECT 15.8000 64.8000 16.2000 65.2000 ;
	    RECT 35.0000 64.8000 35.4000 65.2000 ;
	    RECT 38.2000 65.1000 38.6000 65.2000 ;
	    RECT 43.0000 65.1000 43.4000 65.2000 ;
	    RECT 37.4000 64.8000 43.4000 65.1000 ;
	    RECT 48.6000 65.1000 49.0000 65.2000 ;
	    RECT 57.4000 65.1000 57.8000 65.2000 ;
	    RECT 59.8000 65.1000 60.2000 65.2000 ;
	    RECT 77.4000 65.1000 77.8000 65.2000 ;
	    RECT 87.0000 65.1000 87.4000 65.2000 ;
	    RECT 48.6000 64.8000 63.3000 65.1000 ;
	    RECT 77.4000 64.8000 87.4000 65.1000 ;
	    RECT 96.6000 65.1000 97.0000 65.2000 ;
	    RECT 107.8000 65.1000 108.2000 65.2000 ;
	    RECT 96.6000 64.8000 108.2000 65.1000 ;
	    RECT 109.4000 65.1000 109.7000 65.8000 ;
	    RECT 110.2000 65.1000 110.6000 65.2000 ;
	    RECT 109.4000 64.8000 110.6000 65.1000 ;
	    RECT 115.0000 65.1000 115.4000 65.2000 ;
	    RECT 117.4000 65.1000 117.7000 65.8000 ;
	    RECT 115.0000 64.8000 117.7000 65.1000 ;
	    RECT 118.2000 65.1000 118.6000 65.2000 ;
	    RECT 130.2000 65.1000 130.6000 65.2000 ;
	    RECT 133.4000 65.1000 133.8000 65.2000 ;
	    RECT 139.8000 65.1000 140.2000 65.2000 ;
	    RECT 141.4000 65.1000 141.8000 65.2000 ;
	    RECT 118.2000 64.8000 119.3000 65.1000 ;
	    RECT 130.2000 64.8000 134.5000 65.1000 ;
	    RECT 139.8000 64.8000 141.8000 65.1000 ;
	    RECT 27.0000 64.1000 27.4000 64.2000 ;
	    RECT 33.4000 64.1000 33.8000 64.2000 ;
	    RECT 27.0000 63.8000 33.8000 64.1000 ;
	    RECT 35.0000 64.1000 35.3000 64.8000 ;
	    RECT 63.0000 64.2000 63.3000 64.8000 ;
	    RECT 47.0000 64.1000 47.4000 64.2000 ;
	    RECT 53.4000 64.1000 53.8000 64.2000 ;
	    RECT 55.8000 64.1000 56.2000 64.2000 ;
	    RECT 35.0000 63.8000 56.2000 64.1000 ;
	    RECT 63.0000 63.8000 63.4000 64.2000 ;
	    RECT 106.2000 64.1000 106.6000 64.2000 ;
	    RECT 111.0000 64.1000 111.4000 64.2000 ;
	    RECT 106.2000 63.8000 111.4000 64.1000 ;
	    RECT 116.6000 64.1000 117.0000 64.2000 ;
	    RECT 120.6000 64.1000 121.0000 64.2000 ;
	    RECT 116.6000 63.8000 121.0000 64.1000 ;
	    RECT 94.2000 63.1000 94.6000 63.2000 ;
	    RECT 96.6000 63.1000 97.0000 63.2000 ;
	    RECT 94.2000 62.8000 97.0000 63.1000 ;
	    RECT 107.8000 63.1000 108.2000 63.2000 ;
	    RECT 110.2000 63.1000 110.6000 63.2000 ;
	    RECT 107.8000 62.8000 120.1000 63.1000 ;
	    RECT 119.8000 62.2000 120.1000 62.8000 ;
	    RECT 39.0000 62.1000 39.4000 62.2000 ;
	    RECT 72.6000 62.1000 73.0000 62.2000 ;
	    RECT 39.0000 61.8000 73.0000 62.1000 ;
	    RECT 78.2000 62.1000 78.6000 62.2000 ;
	    RECT 84.6000 62.1000 85.0000 62.2000 ;
	    RECT 78.2000 61.8000 85.0000 62.1000 ;
	    RECT 119.8000 61.8000 120.2000 62.2000 ;
	    RECT 71.8000 61.1000 72.2000 61.2000 ;
	    RECT 78.2000 61.1000 78.6000 61.2000 ;
	    RECT 71.8000 60.8000 78.6000 61.1000 ;
	    RECT 110.2000 61.1000 110.6000 61.2000 ;
	    RECT 121.4000 61.1000 121.8000 61.2000 ;
	    RECT 110.2000 60.8000 121.8000 61.1000 ;
	    RECT 96.6000 60.1000 97.0000 60.2000 ;
	    RECT 103.8000 60.1000 104.2000 60.2000 ;
	    RECT 112.6000 60.1000 113.0000 60.2000 ;
	    RECT 96.6000 59.8000 113.0000 60.1000 ;
	    RECT 6.2000 59.1000 6.6000 59.2000 ;
	    RECT 8.6000 59.1000 9.0000 59.2000 ;
	    RECT 19.0000 59.1000 19.4000 59.2000 ;
	    RECT 6.2000 58.8000 19.4000 59.1000 ;
	    RECT 31.0000 59.1000 31.4000 59.2000 ;
	    RECT 39.8000 59.1000 40.2000 59.2000 ;
	    RECT 31.0000 58.8000 40.2000 59.1000 ;
	    RECT 87.8000 58.8000 88.2000 59.2000 ;
	    RECT 103.0000 59.1000 103.4000 59.2000 ;
	    RECT 121.4000 59.1000 121.8000 59.2000 ;
	    RECT 130.2000 59.1000 130.6000 59.2000 ;
	    RECT 103.0000 58.8000 119.3000 59.1000 ;
	    RECT 121.4000 58.8000 130.6000 59.1000 ;
	    RECT 29.4000 58.1000 29.8000 58.2000 ;
	    RECT 34.2000 58.1000 34.6000 58.2000 ;
	    RECT 54.2000 58.1000 54.6000 58.2000 ;
	    RECT 29.4000 57.8000 54.6000 58.1000 ;
	    RECT 87.8000 58.1000 88.1000 58.8000 ;
	    RECT 119.0000 58.2000 119.3000 58.8000 ;
	    RECT 91.8000 58.1000 92.2000 58.2000 ;
	    RECT 87.8000 57.8000 92.2000 58.1000 ;
	    RECT 113.4000 57.8000 113.8000 58.2000 ;
	    RECT 119.0000 57.8000 119.4000 58.2000 ;
	    RECT 123.8000 58.1000 124.2000 58.2000 ;
	    RECT 124.6000 58.1000 125.0000 58.2000 ;
	    RECT 123.8000 57.8000 125.0000 58.1000 ;
	    RECT 125.4000 57.8000 125.8000 58.2000 ;
	    RECT 58.2000 56.8000 58.6000 57.2000 ;
	    RECT 84.6000 57.1000 85.0000 57.2000 ;
	    RECT 94.2000 57.1000 94.6000 57.2000 ;
	    RECT 84.6000 56.8000 94.6000 57.1000 ;
	    RECT 113.4000 57.1000 113.7000 57.8000 ;
	    RECT 119.0000 57.1000 119.4000 57.2000 ;
	    RECT 113.4000 56.8000 119.4000 57.1000 ;
	    RECT 123.0000 57.1000 123.4000 57.2000 ;
	    RECT 125.4000 57.1000 125.7000 57.8000 ;
	    RECT 123.0000 56.8000 125.7000 57.1000 ;
	    RECT 15.8000 55.8000 16.2000 56.2000 ;
	    RECT 23.8000 56.1000 24.2000 56.2000 ;
	    RECT 41.4000 56.1000 41.8000 56.2000 ;
	    RECT 58.2000 56.1000 58.5000 56.8000 ;
	    RECT 23.8000 55.8000 58.5000 56.1000 ;
	    RECT 90.2000 56.1000 90.6000 56.2000 ;
	    RECT 91.0000 56.1000 91.4000 56.2000 ;
	    RECT 90.2000 55.8000 91.4000 56.1000 ;
	    RECT 92.6000 56.1000 93.0000 56.2000 ;
	    RECT 101.4000 56.1000 101.8000 56.2000 ;
	    RECT 92.6000 55.8000 101.8000 56.1000 ;
	    RECT 113.4000 56.1000 113.8000 56.2000 ;
	    RECT 114.2000 56.1000 114.6000 56.2000 ;
	    RECT 113.4000 55.8000 114.6000 56.1000 ;
	    RECT 123.8000 56.1000 124.2000 56.2000 ;
	    RECT 130.2000 56.1000 130.6000 56.2000 ;
	    RECT 123.8000 55.8000 130.6000 56.1000 ;
	    RECT 5.4000 55.1000 5.8000 55.2000 ;
	    RECT 9.4000 55.1000 9.8000 55.2000 ;
	    RECT 12.6000 55.1000 13.0000 55.2000 ;
	    RECT 5.4000 54.8000 13.0000 55.1000 ;
	    RECT 15.8000 55.1000 16.1000 55.8000 ;
	    RECT 21.4000 55.1000 21.8000 55.2000 ;
	    RECT 15.8000 54.8000 21.8000 55.1000 ;
	    RECT 35.0000 55.1000 35.4000 55.2000 ;
	    RECT 36.6000 55.1000 37.0000 55.2000 ;
	    RECT 35.0000 54.8000 37.0000 55.1000 ;
	    RECT 42.2000 54.8000 42.6000 55.2000 ;
	    RECT 43.8000 55.1000 44.2000 55.2000 ;
	    RECT 47.0000 55.1000 47.4000 55.2000 ;
	    RECT 43.8000 54.8000 47.4000 55.1000 ;
	    RECT 55.0000 55.1000 55.4000 55.2000 ;
	    RECT 64.6000 55.1000 65.0000 55.2000 ;
	    RECT 69.4000 55.1000 69.8000 55.2000 ;
	    RECT 55.0000 54.8000 69.8000 55.1000 ;
	    RECT 71.0000 55.1000 71.4000 55.2000 ;
	    RECT 82.2000 55.1000 82.6000 55.2000 ;
	    RECT 71.0000 54.8000 82.6000 55.1000 ;
	    RECT 86.2000 55.1000 86.6000 55.2000 ;
	    RECT 90.2000 55.1000 90.6000 55.2000 ;
	    RECT 86.2000 54.8000 90.6000 55.1000 ;
	    RECT 113.4000 55.1000 113.8000 55.2000 ;
	    RECT 115.0000 55.1000 115.4000 55.2000 ;
	    RECT 124.6000 55.1000 125.0000 55.2000 ;
	    RECT 113.4000 54.8000 125.0000 55.1000 ;
	    RECT 127.8000 55.1000 128.2000 55.2000 ;
	    RECT 138.2000 55.1000 138.6000 55.2000 ;
	    RECT 140.6000 55.1000 141.0000 55.2000 ;
	    RECT 144.6000 55.1000 145.0000 55.2000 ;
	    RECT 145.4000 55.1000 145.8000 55.2000 ;
	    RECT 127.8000 54.8000 145.8000 55.1000 ;
	    RECT 17.4000 54.1000 17.8000 54.2000 ;
	    RECT 40.6000 54.1000 41.0000 54.2000 ;
	    RECT 42.2000 54.1000 42.5000 54.8000 ;
	    RECT 17.4000 53.8000 25.7000 54.1000 ;
	    RECT 40.6000 53.8000 42.5000 54.1000 ;
	    RECT 43.0000 54.1000 43.4000 54.2000 ;
	    RECT 54.2000 54.1000 54.6000 54.2000 ;
	    RECT 43.0000 53.8000 54.6000 54.1000 ;
	    RECT 60.6000 54.1000 61.0000 54.2000 ;
	    RECT 63.8000 54.1000 64.2000 54.2000 ;
	    RECT 60.6000 53.8000 64.2000 54.1000 ;
	    RECT 68.6000 54.1000 69.0000 54.2000 ;
	    RECT 70.2000 54.1000 70.6000 54.2000 ;
	    RECT 68.6000 53.8000 70.6000 54.1000 ;
	    RECT 75.8000 54.1000 76.2000 54.2000 ;
	    RECT 125.4000 54.1000 125.8000 54.2000 ;
	    RECT 127.0000 54.1000 127.4000 54.2000 ;
	    RECT 75.8000 53.8000 127.4000 54.1000 ;
	    RECT 131.8000 54.1000 132.2000 54.2000 ;
	    RECT 143.8000 54.1000 144.2000 54.2000 ;
	    RECT 131.8000 53.8000 144.2000 54.1000 ;
	    RECT 25.4000 53.2000 25.7000 53.8000 ;
	    RECT 0.6000 53.1000 1.0000 53.2000 ;
	    RECT 2.2000 53.1000 2.6000 53.2000 ;
	    RECT 4.6000 53.1000 5.0000 53.2000 ;
	    RECT 0.6000 52.8000 5.0000 53.1000 ;
	    RECT 25.4000 52.8000 25.8000 53.2000 ;
	    RECT 39.8000 53.1000 40.2000 53.2000 ;
	    RECT 49.4000 53.1000 49.8000 53.2000 ;
	    RECT 39.8000 52.8000 49.8000 53.1000 ;
	    RECT 65.4000 53.1000 65.8000 53.2000 ;
	    RECT 74.2000 53.1000 74.6000 53.2000 ;
	    RECT 65.4000 52.8000 74.6000 53.1000 ;
	    RECT 76.6000 53.1000 77.0000 53.2000 ;
	    RECT 91.0000 53.1000 91.4000 53.2000 ;
	    RECT 76.6000 52.8000 91.4000 53.1000 ;
	    RECT 92.6000 53.1000 93.0000 53.2000 ;
	    RECT 93.4000 53.1000 93.8000 53.2000 ;
	    RECT 92.6000 52.8000 93.8000 53.1000 ;
	    RECT 100.6000 53.1000 101.0000 53.2000 ;
	    RECT 111.8000 53.1000 112.2000 53.2000 ;
	    RECT 124.6000 53.1000 125.0000 53.2000 ;
	    RECT 131.8000 53.1000 132.2000 53.2000 ;
	    RECT 100.6000 52.8000 132.2000 53.1000 ;
	    RECT 143.0000 53.1000 143.4000 53.2000 ;
	    RECT 145.4000 53.1000 145.8000 53.2000 ;
	    RECT 143.0000 52.8000 145.8000 53.1000 ;
	    RECT 23.0000 52.1000 23.4000 52.2000 ;
	    RECT 27.0000 52.1000 27.4000 52.2000 ;
	    RECT 23.0000 51.8000 27.4000 52.1000 ;
	    RECT 30.2000 52.1000 30.6000 52.2000 ;
	    RECT 63.0000 52.1000 63.4000 52.2000 ;
	    RECT 71.8000 52.1000 72.2000 52.2000 ;
	    RECT 72.6000 52.1000 73.0000 52.2000 ;
	    RECT 77.4000 52.1000 77.8000 52.2000 ;
	    RECT 30.2000 51.8000 77.8000 52.1000 ;
	    RECT 79.8000 52.1000 80.2000 52.2000 ;
	    RECT 81.4000 52.1000 81.8000 52.2000 ;
	    RECT 79.8000 51.8000 81.8000 52.1000 ;
	    RECT 82.2000 52.1000 82.6000 52.2000 ;
	    RECT 87.0000 52.1000 87.4000 52.2000 ;
	    RECT 82.2000 51.8000 87.4000 52.1000 ;
	    RECT 89.4000 52.1000 89.8000 52.2000 ;
	    RECT 90.2000 52.1000 90.6000 52.2000 ;
	    RECT 108.6000 52.1000 109.0000 52.2000 ;
	    RECT 114.2000 52.1000 114.6000 52.2000 ;
	    RECT 89.4000 51.8000 90.6000 52.1000 ;
	    RECT 91.0000 51.8000 114.6000 52.1000 ;
	    RECT 36.6000 51.1000 37.0000 51.2000 ;
	    RECT 42.2000 51.1000 42.6000 51.2000 ;
	    RECT 36.6000 50.8000 42.6000 51.1000 ;
	    RECT 83.0000 51.1000 83.4000 51.2000 ;
	    RECT 91.0000 51.1000 91.3000 51.8000 ;
	    RECT 83.0000 50.8000 91.3000 51.1000 ;
	    RECT 102.2000 51.1000 102.6000 51.2000 ;
	    RECT 130.2000 51.1000 130.6000 51.2000 ;
	    RECT 134.2000 51.1000 134.6000 51.2000 ;
	    RECT 135.8000 51.1000 136.2000 51.2000 ;
	    RECT 102.2000 50.8000 136.2000 51.1000 ;
	    RECT 18.2000 50.1000 18.6000 50.2000 ;
	    RECT 25.4000 50.1000 25.8000 50.2000 ;
	    RECT 31.0000 50.1000 31.4000 50.2000 ;
	    RECT 64.6000 50.1000 65.0000 50.2000 ;
	    RECT 69.4000 50.1000 69.8000 50.2000 ;
	    RECT 18.2000 49.8000 69.8000 50.1000 ;
	    RECT 80.6000 50.1000 81.0000 50.2000 ;
	    RECT 83.0000 50.1000 83.4000 50.2000 ;
	    RECT 80.6000 49.8000 83.4000 50.1000 ;
	    RECT 83.8000 50.1000 84.2000 50.2000 ;
	    RECT 89.4000 50.1000 89.8000 50.2000 ;
	    RECT 83.8000 49.8000 89.8000 50.1000 ;
	    RECT 133.4000 50.1000 133.8000 50.2000 ;
	    RECT 142.2000 50.1000 142.6000 50.2000 ;
	    RECT 133.4000 49.8000 142.6000 50.1000 ;
	    RECT 6.2000 49.1000 6.6000 49.2000 ;
	    RECT 10.2000 49.1000 10.6000 49.2000 ;
	    RECT 6.2000 48.8000 10.6000 49.1000 ;
	    RECT 73.4000 48.8000 73.8000 49.2000 ;
	    RECT 79.0000 49.1000 79.4000 49.2000 ;
	    RECT 82.2000 49.1000 82.6000 49.2000 ;
	    RECT 79.0000 48.8000 82.6000 49.1000 ;
	    RECT 83.8000 49.1000 84.2000 49.2000 ;
	    RECT 91.0000 49.1000 91.4000 49.2000 ;
	    RECT 83.8000 48.8000 91.4000 49.1000 ;
	    RECT 93.4000 49.1000 93.8000 49.2000 ;
	    RECT 94.2000 49.1000 94.6000 49.2000 ;
	    RECT 93.4000 48.8000 94.6000 49.1000 ;
	    RECT 127.0000 49.1000 127.4000 49.2000 ;
	    RECT 130.2000 49.1000 130.6000 49.2000 ;
	    RECT 140.6000 49.1000 141.0000 49.2000 ;
	    RECT 127.0000 48.8000 141.0000 49.1000 ;
	    RECT 8.6000 48.1000 9.0000 48.2000 ;
	    RECT 17.4000 48.1000 17.8000 48.2000 ;
	    RECT 8.6000 47.8000 17.8000 48.1000 ;
	    RECT 24.6000 48.1000 25.0000 48.2000 ;
	    RECT 28.6000 48.1000 29.0000 48.2000 ;
	    RECT 61.4000 48.1000 61.8000 48.2000 ;
	    RECT 63.0000 48.1000 63.4000 48.2000 ;
	    RECT 65.4000 48.1000 65.8000 48.2000 ;
	    RECT 67.0000 48.1000 67.4000 48.2000 ;
	    RECT 24.6000 47.8000 67.4000 48.1000 ;
	    RECT 71.0000 48.1000 71.4000 48.2000 ;
	    RECT 73.4000 48.1000 73.7000 48.8000 ;
	    RECT 71.0000 47.8000 73.7000 48.1000 ;
	    RECT 75.8000 48.1000 76.2000 48.2000 ;
	    RECT 101.4000 48.1000 101.8000 48.2000 ;
	    RECT 75.8000 47.8000 101.8000 48.1000 ;
	    RECT 120.6000 48.1000 121.0000 48.2000 ;
	    RECT 135.8000 48.1000 136.2000 48.2000 ;
	    RECT 120.6000 47.8000 136.2000 48.1000 ;
	    RECT 7.0000 47.1000 7.4000 47.2000 ;
	    RECT 10.2000 47.1000 10.6000 47.2000 ;
	    RECT 7.0000 46.8000 10.6000 47.1000 ;
	    RECT 11.8000 47.1000 12.2000 47.2000 ;
	    RECT 15.0000 47.1000 15.4000 47.2000 ;
	    RECT 15.8000 47.1000 16.2000 47.2000 ;
	    RECT 11.8000 46.8000 16.2000 47.1000 ;
	    RECT 20.6000 47.1000 21.0000 47.2000 ;
	    RECT 34.2000 47.1000 34.6000 47.2000 ;
	    RECT 20.6000 46.8000 34.6000 47.1000 ;
	    RECT 64.6000 47.1000 65.0000 47.2000 ;
	    RECT 75.0000 47.1000 75.4000 47.2000 ;
	    RECT 64.6000 46.8000 75.4000 47.1000 ;
	    RECT 75.8000 46.8000 76.2000 47.2000 ;
	    RECT 90.2000 46.8000 90.6000 47.2000 ;
	    RECT 91.0000 47.1000 91.4000 47.2000 ;
	    RECT 96.6000 47.1000 97.0000 47.2000 ;
	    RECT 91.0000 46.8000 97.0000 47.1000 ;
	    RECT 107.8000 47.1000 108.2000 47.2000 ;
	    RECT 121.4000 47.1000 121.8000 47.2000 ;
	    RECT 129.4000 47.1000 129.8000 47.2000 ;
	    RECT 107.8000 46.8000 118.5000 47.1000 ;
	    RECT 121.4000 46.8000 129.8000 47.1000 ;
	    RECT 135.8000 47.1000 136.2000 47.2000 ;
	    RECT 139.8000 47.1000 140.2000 47.2000 ;
	    RECT 135.8000 46.8000 140.2000 47.1000 ;
	    RECT 25.4000 46.1000 25.8000 46.2000 ;
	    RECT 33.4000 46.1000 33.8000 46.2000 ;
	    RECT 44.6000 46.1000 45.0000 46.2000 ;
	    RECT 25.4000 45.8000 33.8000 46.1000 ;
	    RECT 43.0000 45.8000 45.0000 46.1000 ;
	    RECT 68.6000 45.8000 69.0000 46.2000 ;
	    RECT 73.4000 46.1000 73.8000 46.2000 ;
	    RECT 75.8000 46.1000 76.1000 46.8000 ;
	    RECT 73.4000 45.8000 76.1000 46.1000 ;
	    RECT 86.2000 46.1000 86.6000 46.2000 ;
	    RECT 90.2000 46.1000 90.5000 46.8000 ;
	    RECT 118.2000 46.2000 118.5000 46.8000 ;
	    RECT 86.2000 45.8000 90.5000 46.1000 ;
	    RECT 91.0000 46.1000 91.4000 46.2000 ;
	    RECT 99.8000 46.1000 100.2000 46.2000 ;
	    RECT 91.0000 45.8000 100.2000 46.1000 ;
	    RECT 118.2000 45.8000 118.6000 46.2000 ;
	    RECT 124.6000 46.1000 125.0000 46.2000 ;
	    RECT 126.2000 46.1000 126.6000 46.2000 ;
	    RECT 124.6000 45.8000 126.6000 46.1000 ;
	    RECT 127.8000 46.1000 128.2000 46.2000 ;
	    RECT 131.0000 46.1000 131.4000 46.2000 ;
	    RECT 127.8000 45.8000 131.4000 46.1000 ;
	    RECT 43.0000 45.2000 43.3000 45.8000 ;
	    RECT 12.6000 45.1000 13.0000 45.2000 ;
	    RECT 16.6000 45.1000 17.0000 45.2000 ;
	    RECT 20.6000 45.1000 21.0000 45.2000 ;
	    RECT 12.6000 44.8000 21.0000 45.1000 ;
	    RECT 27.8000 44.8000 28.2000 45.2000 ;
	    RECT 43.0000 44.8000 43.4000 45.2000 ;
	    RECT 56.6000 45.1000 57.0000 45.2000 ;
	    RECT 63.8000 45.1000 64.2000 45.2000 ;
	    RECT 45.4000 44.8000 64.2000 45.1000 ;
	    RECT 68.6000 45.1000 68.9000 45.8000 ;
	    RECT 77.4000 45.1000 77.8000 45.2000 ;
	    RECT 68.6000 44.8000 77.8000 45.1000 ;
	    RECT 79.8000 45.1000 80.2000 45.2000 ;
	    RECT 83.8000 45.1000 84.2000 45.2000 ;
	    RECT 89.4000 45.1000 89.8000 45.2000 ;
	    RECT 79.8000 44.8000 89.8000 45.1000 ;
	    RECT 95.0000 45.1000 95.4000 45.2000 ;
	    RECT 95.8000 45.1000 96.2000 45.2000 ;
	    RECT 95.0000 44.8000 96.2000 45.1000 ;
	    RECT 140.6000 45.1000 141.0000 45.2000 ;
	    RECT 141.4000 45.1000 141.8000 45.2000 ;
	    RECT 140.6000 44.8000 141.8000 45.1000 ;
	    RECT 19.0000 44.1000 19.4000 44.2000 ;
	    RECT 26.2000 44.1000 26.6000 44.2000 ;
	    RECT 27.8000 44.1000 28.1000 44.8000 ;
	    RECT 19.0000 43.8000 28.1000 44.1000 ;
	    RECT 29.4000 44.1000 29.8000 44.2000 ;
	    RECT 34.2000 44.1000 34.6000 44.2000 ;
	    RECT 45.4000 44.1000 45.7000 44.8000 ;
	    RECT 29.4000 43.8000 45.7000 44.1000 ;
	    RECT 57.4000 44.1000 57.8000 44.2000 ;
	    RECT 59.8000 44.1000 60.2000 44.2000 ;
	    RECT 57.4000 43.8000 60.2000 44.1000 ;
	    RECT 74.2000 44.1000 74.6000 44.2000 ;
	    RECT 81.4000 44.1000 81.8000 44.2000 ;
	    RECT 91.8000 44.1000 92.2000 44.2000 ;
	    RECT 94.2000 44.1000 94.6000 44.2000 ;
	    RECT 108.6000 44.1000 109.0000 44.2000 ;
	    RECT 74.2000 43.8000 81.8000 44.1000 ;
	    RECT 88.6000 43.8000 92.2000 44.1000 ;
	    RECT 92.6000 43.8000 94.6000 44.1000 ;
	    RECT 95.8000 43.8000 109.0000 44.1000 ;
	    RECT 138.2000 44.1000 138.6000 44.2000 ;
	    RECT 139.8000 44.1000 140.2000 44.2000 ;
	    RECT 138.2000 43.8000 140.2000 44.1000 ;
	    RECT 88.6000 43.2000 88.9000 43.8000 ;
	    RECT 92.6000 43.2000 92.9000 43.8000 ;
	    RECT 95.8000 43.2000 96.1000 43.8000 ;
	    RECT 88.6000 42.8000 89.0000 43.2000 ;
	    RECT 92.6000 42.8000 93.0000 43.2000 ;
	    RECT 95.8000 42.8000 96.2000 43.2000 ;
	    RECT 53.4000 42.1000 53.8000 42.2000 ;
	    RECT 94.2000 42.1000 94.6000 42.2000 ;
	    RECT 53.4000 41.8000 94.6000 42.1000 ;
	    RECT 103.0000 41.2000 103.3000 42.1000 ;
	    RECT 103.0000 40.8000 103.4000 41.2000 ;
	    RECT 35.8000 39.1000 36.2000 39.2000 ;
	    RECT 52.6000 39.1000 53.0000 39.2000 ;
	    RECT 35.8000 38.8000 53.0000 39.1000 ;
	    RECT 55.0000 39.1000 55.4000 39.2000 ;
	    RECT 76.6000 39.1000 77.0000 39.2000 ;
	    RECT 55.0000 38.8000 77.0000 39.1000 ;
	    RECT 77.4000 39.1000 77.8000 39.2000 ;
	    RECT 91.0000 39.1000 91.4000 39.2000 ;
	    RECT 77.4000 38.8000 91.4000 39.1000 ;
	    RECT 109.4000 39.1000 109.8000 39.2000 ;
	    RECT 121.4000 39.1000 121.8000 39.2000 ;
	    RECT 109.4000 38.8000 121.8000 39.1000 ;
	    RECT 13.4000 38.1000 13.8000 38.2000 ;
	    RECT 23.8000 38.1000 24.2000 38.2000 ;
	    RECT 13.4000 37.8000 24.2000 38.1000 ;
	    RECT 34.2000 38.1000 34.6000 38.2000 ;
	    RECT 58.2000 38.1000 58.6000 38.2000 ;
	    RECT 34.2000 37.8000 58.6000 38.1000 ;
	    RECT 63.0000 38.1000 63.4000 38.2000 ;
	    RECT 67.0000 38.1000 67.4000 38.2000 ;
	    RECT 79.8000 38.1000 80.2000 38.2000 ;
	    RECT 63.0000 37.8000 80.2000 38.1000 ;
	    RECT 100.6000 38.1000 101.0000 38.2000 ;
	    RECT 105.4000 38.1000 105.8000 38.2000 ;
	    RECT 100.6000 37.8000 105.8000 38.1000 ;
	    RECT 106.2000 38.1000 106.6000 38.2000 ;
	    RECT 120.6000 38.1000 121.0000 38.2000 ;
	    RECT 106.2000 37.8000 121.0000 38.1000 ;
	    RECT 23.0000 37.1000 23.4000 37.2000 ;
	    RECT 23.0000 36.8000 25.7000 37.1000 ;
	    RECT 25.4000 36.2000 25.7000 36.8000 ;
	    RECT 40.6000 36.8000 41.0000 37.2000 ;
	    RECT 72.6000 37.1000 73.0000 37.2000 ;
	    RECT 75.0000 37.1000 75.4000 37.2000 ;
	    RECT 72.6000 36.8000 75.4000 37.1000 ;
	    RECT 77.4000 37.1000 77.8000 37.2000 ;
	    RECT 79.0000 37.1000 79.4000 37.2000 ;
	    RECT 77.4000 36.8000 79.4000 37.1000 ;
	    RECT 79.8000 37.1000 80.2000 37.2000 ;
	    RECT 83.0000 37.1000 83.4000 37.2000 ;
	    RECT 107.0000 37.1000 107.4000 37.2000 ;
	    RECT 79.8000 36.8000 107.4000 37.1000 ;
	    RECT 111.0000 37.1000 111.4000 37.2000 ;
	    RECT 134.2000 37.1000 134.6000 37.2000 ;
	    RECT 111.0000 36.8000 134.6000 37.1000 ;
	    RECT 9.4000 35.8000 9.8000 36.2000 ;
	    RECT 25.4000 35.8000 25.8000 36.2000 ;
	    RECT 27.8000 35.8000 28.2000 36.2000 ;
	    RECT 32.6000 36.1000 33.0000 36.2000 ;
	    RECT 37.4000 36.1000 37.8000 36.2000 ;
	    RECT 40.6000 36.1000 40.9000 36.8000 ;
	    RECT 32.6000 35.8000 40.9000 36.1000 ;
	    RECT 51.8000 36.1000 52.2000 36.2000 ;
	    RECT 84.6000 36.1000 85.0000 36.2000 ;
	    RECT 51.8000 35.8000 85.0000 36.1000 ;
	    RECT 89.4000 36.1000 89.8000 36.2000 ;
	    RECT 102.2000 36.1000 102.6000 36.2000 ;
	    RECT 104.6000 36.1000 105.0000 36.2000 ;
	    RECT 109.4000 36.1000 109.8000 36.2000 ;
	    RECT 89.4000 35.8000 102.6000 36.1000 ;
	    RECT 103.8000 35.8000 109.8000 36.1000 ;
	    RECT 110.2000 36.1000 110.6000 36.2000 ;
	    RECT 114.2000 36.1000 114.6000 36.2000 ;
	    RECT 110.2000 35.8000 114.6000 36.1000 ;
	    RECT 115.8000 36.1000 116.2000 36.2000 ;
	    RECT 122.2000 36.1000 122.6000 36.2000 ;
	    RECT 127.8000 36.1000 128.2000 36.2000 ;
	    RECT 135.0000 36.1000 135.4000 36.2000 ;
	    RECT 137.4000 36.1000 137.8000 36.2000 ;
	    RECT 115.8000 35.8000 137.8000 36.1000 ;
	    RECT 9.4000 35.1000 9.7000 35.8000 ;
	    RECT 14.2000 35.1000 14.6000 35.2000 ;
	    RECT 9.4000 34.8000 14.6000 35.1000 ;
	    RECT 19.8000 35.1000 20.2000 35.2000 ;
	    RECT 22.2000 35.1000 22.6000 35.2000 ;
	    RECT 19.8000 34.8000 22.6000 35.1000 ;
	    RECT 27.0000 35.1000 27.4000 35.2000 ;
	    RECT 27.8000 35.1000 28.1000 35.8000 ;
	    RECT 27.0000 34.8000 28.1000 35.1000 ;
	    RECT 28.6000 35.1000 29.0000 35.2000 ;
	    RECT 34.2000 35.1000 34.6000 35.2000 ;
	    RECT 28.6000 34.8000 34.6000 35.1000 ;
	    RECT 39.8000 35.1000 40.2000 35.2000 ;
	    RECT 46.2000 35.1000 46.6000 35.2000 ;
	    RECT 39.8000 34.8000 46.6000 35.1000 ;
	    RECT 47.8000 35.1000 48.2000 35.2000 ;
	    RECT 53.4000 35.1000 53.8000 35.2000 ;
	    RECT 47.8000 34.8000 53.8000 35.1000 ;
	    RECT 58.2000 35.1000 58.6000 35.2000 ;
	    RECT 60.6000 35.1000 61.0000 35.2000 ;
	    RECT 58.2000 34.8000 61.0000 35.1000 ;
	    RECT 69.4000 35.1000 69.8000 35.2000 ;
	    RECT 74.2000 35.1000 74.6000 35.2000 ;
	    RECT 76.6000 35.1000 77.0000 35.2000 ;
	    RECT 69.4000 34.8000 77.0000 35.1000 ;
	    RECT 78.2000 35.1000 78.6000 35.2000 ;
	    RECT 89.4000 35.1000 89.8000 35.2000 ;
	    RECT 78.2000 34.8000 89.8000 35.1000 ;
	    RECT 103.8000 35.1000 104.2000 35.2000 ;
	    RECT 106.2000 35.1000 106.6000 35.2000 ;
	    RECT 103.8000 34.8000 106.6000 35.1000 ;
	    RECT 112.6000 34.8000 113.0000 35.2000 ;
	    RECT 125.4000 34.8000 125.8000 35.2000 ;
	    RECT 128.6000 35.1000 129.0000 35.2000 ;
	    RECT 131.8000 35.1000 132.2000 35.2000 ;
	    RECT 128.6000 34.8000 132.2000 35.1000 ;
	    RECT 133.4000 35.1000 133.8000 35.2000 ;
	    RECT 136.6000 35.1000 137.0000 35.2000 ;
	    RECT 133.4000 34.8000 137.0000 35.1000 ;
	    RECT 140.6000 34.8000 141.0000 35.2000 ;
	    RECT 6.2000 33.8000 6.6000 34.2000 ;
	    RECT 12.6000 33.8000 13.0000 34.2000 ;
	    RECT 17.4000 34.1000 17.8000 34.2000 ;
	    RECT 21.4000 34.1000 21.8000 34.2000 ;
	    RECT 30.2000 34.1000 30.6000 34.2000 ;
	    RECT 17.4000 33.8000 30.6000 34.1000 ;
	    RECT 63.8000 34.1000 64.2000 34.2000 ;
	    RECT 75.8000 34.1000 76.2000 34.2000 ;
	    RECT 87.8000 34.1000 88.2000 34.2000 ;
	    RECT 63.8000 33.8000 88.2000 34.1000 ;
	    RECT 99.8000 34.1000 100.2000 34.2000 ;
	    RECT 107.0000 34.1000 107.4000 34.2000 ;
	    RECT 112.6000 34.1000 112.9000 34.8000 ;
	    RECT 125.4000 34.1000 125.7000 34.8000 ;
	    RECT 140.6000 34.2000 140.9000 34.8000 ;
	    RECT 136.6000 34.1000 137.0000 34.2000 ;
	    RECT 99.8000 33.8000 137.0000 34.1000 ;
	    RECT 140.6000 33.8000 141.0000 34.2000 ;
	    RECT 6.2000 33.1000 6.5000 33.8000 ;
	    RECT 12.6000 33.1000 12.9000 33.8000 ;
	    RECT 6.2000 32.8000 12.9000 33.1000 ;
	    RECT 28.6000 33.1000 29.0000 33.2000 ;
	    RECT 32.6000 33.1000 33.0000 33.2000 ;
	    RECT 28.6000 32.8000 33.0000 33.1000 ;
	    RECT 45.4000 33.1000 45.8000 33.2000 ;
	    RECT 51.8000 33.1000 52.2000 33.2000 ;
	    RECT 57.4000 33.1000 57.8000 33.2000 ;
	    RECT 45.4000 32.8000 57.8000 33.1000 ;
	    RECT 59.8000 33.1000 60.2000 33.2000 ;
	    RECT 66.2000 33.1000 66.6000 33.2000 ;
	    RECT 59.8000 32.8000 66.6000 33.1000 ;
	    RECT 67.8000 33.1000 68.2000 33.2000 ;
	    RECT 68.6000 33.1000 69.0000 33.2000 ;
	    RECT 71.0000 33.1000 71.4000 33.2000 ;
	    RECT 67.8000 32.8000 71.4000 33.1000 ;
	    RECT 86.2000 33.1000 86.6000 33.2000 ;
	    RECT 87.8000 33.1000 88.2000 33.2000 ;
	    RECT 86.2000 32.8000 88.2000 33.1000 ;
	    RECT 102.2000 33.1000 102.6000 33.2000 ;
	    RECT 105.4000 33.1000 105.8000 33.2000 ;
	    RECT 128.6000 33.1000 129.0000 33.2000 ;
	    RECT 102.2000 32.8000 105.8000 33.1000 ;
	    RECT 123.8000 32.8000 129.0000 33.1000 ;
	    RECT 139.8000 33.1000 140.2000 33.2000 ;
	    RECT 141.4000 33.1000 141.8000 33.2000 ;
	    RECT 144.6000 33.1000 145.0000 33.2000 ;
	    RECT 139.8000 32.8000 145.0000 33.1000 ;
	    RECT 123.8000 32.2000 124.1000 32.8000 ;
	    RECT 17.4000 32.1000 17.8000 32.2000 ;
	    RECT 42.2000 32.1000 42.6000 32.2000 ;
	    RECT 17.4000 31.8000 42.6000 32.1000 ;
	    RECT 43.0000 32.1000 43.4000 32.2000 ;
	    RECT 59.8000 32.1000 60.2000 32.2000 ;
	    RECT 43.0000 31.8000 60.2000 32.1000 ;
	    RECT 60.6000 32.1000 61.0000 32.2000 ;
	    RECT 67.8000 32.1000 68.2000 32.2000 ;
	    RECT 60.6000 31.8000 68.2000 32.1000 ;
	    RECT 123.8000 31.8000 124.2000 32.2000 ;
	    RECT 143.8000 32.1000 144.2000 32.2000 ;
	    RECT 146.2000 32.1000 146.6000 32.2000 ;
	    RECT 143.8000 31.8000 146.6000 32.1000 ;
	    RECT 31.0000 31.1000 31.4000 31.2000 ;
	    RECT 37.4000 31.1000 37.8000 31.2000 ;
	    RECT 31.0000 30.8000 37.8000 31.1000 ;
	    RECT 46.2000 31.1000 46.6000 31.2000 ;
	    RECT 53.4000 31.1000 53.8000 31.2000 ;
	    RECT 69.4000 31.1000 69.8000 31.2000 ;
	    RECT 46.2000 30.8000 69.8000 31.1000 ;
	    RECT 0.6000 30.1000 1.0000 30.2000 ;
	    RECT 24.6000 30.1000 25.0000 30.2000 ;
	    RECT 0.6000 29.8000 25.0000 30.1000 ;
	    RECT 31.8000 30.1000 32.2000 30.2000 ;
	    RECT 46.2000 30.1000 46.6000 30.2000 ;
	    RECT 31.8000 29.8000 46.6000 30.1000 ;
	    RECT 51.8000 30.1000 52.2000 30.2000 ;
	    RECT 72.6000 30.1000 73.0000 30.2000 ;
	    RECT 51.8000 29.8000 73.0000 30.1000 ;
	    RECT 20.6000 29.1000 21.0000 29.2000 ;
	    RECT 27.0000 29.1000 27.4000 29.2000 ;
	    RECT 20.6000 28.8000 27.4000 29.1000 ;
	    RECT 63.8000 29.1000 64.2000 29.2000 ;
	    RECT 81.4000 29.1000 81.8000 29.2000 ;
	    RECT 63.8000 28.8000 81.8000 29.1000 ;
	    RECT 93.4000 29.1000 93.8000 29.2000 ;
	    RECT 98.2000 29.1000 98.6000 29.2000 ;
	    RECT 93.4000 28.8000 98.6000 29.1000 ;
	    RECT 133.4000 29.1000 133.8000 29.2000 ;
	    RECT 135.0000 29.1000 135.4000 29.2000 ;
	    RECT 133.4000 28.8000 135.4000 29.1000 ;
	    RECT 135.8000 29.1000 136.2000 29.2000 ;
	    RECT 139.0000 29.1000 139.4000 29.2000 ;
	    RECT 135.8000 28.8000 139.4000 29.1000 ;
	    RECT 19.8000 28.1000 20.2000 28.2000 ;
	    RECT 41.4000 28.1000 41.8000 28.2000 ;
	    RECT 19.8000 27.8000 41.8000 28.1000 ;
	    RECT 43.8000 28.1000 44.2000 28.2000 ;
	    RECT 51.0000 28.1000 51.4000 28.2000 ;
	    RECT 51.8000 28.1000 52.2000 28.2000 ;
	    RECT 43.8000 27.8000 52.2000 28.1000 ;
	    RECT 54.2000 28.1000 54.6000 28.2000 ;
	    RECT 59.8000 28.1000 60.2000 28.2000 ;
	    RECT 54.2000 27.8000 60.2000 28.1000 ;
	    RECT 65.4000 28.1000 65.8000 28.2000 ;
	    RECT 75.8000 28.1000 76.2000 28.2000 ;
	    RECT 65.4000 27.8000 76.2000 28.1000 ;
	    RECT 76.6000 28.1000 77.0000 28.2000 ;
	    RECT 79.8000 28.1000 80.2000 28.2000 ;
	    RECT 96.6000 28.1000 97.0000 28.2000 ;
	    RECT 76.6000 27.8000 97.0000 28.1000 ;
	    RECT 119.0000 27.8000 119.4000 28.2000 ;
	    RECT 127.0000 28.1000 127.4000 28.2000 ;
	    RECT 130.2000 28.1000 130.6000 28.2000 ;
	    RECT 145.4000 28.1000 145.8000 28.2000 ;
	    RECT 127.0000 27.8000 145.8000 28.1000 ;
	    RECT 7.0000 26.8000 7.4000 27.2000 ;
	    RECT 19.8000 27.1000 20.2000 27.2000 ;
	    RECT 19.8000 26.8000 20.9000 27.1000 ;
	    RECT 7.0000 26.1000 7.3000 26.8000 ;
	    RECT 20.6000 26.2000 20.9000 26.8000 ;
	    RECT 31.0000 26.8000 31.4000 27.2000 ;
	    RECT 35.8000 27.1000 36.2000 27.2000 ;
	    RECT 38.2000 27.1000 38.6000 27.2000 ;
	    RECT 35.8000 26.8000 38.6000 27.1000 ;
	    RECT 42.2000 27.1000 42.6000 27.2000 ;
	    RECT 44.6000 27.1000 45.0000 27.2000 ;
	    RECT 42.2000 26.8000 45.0000 27.1000 ;
	    RECT 45.4000 27.1000 45.8000 27.2000 ;
	    RECT 54.2000 27.1000 54.6000 27.2000 ;
	    RECT 45.4000 26.8000 54.6000 27.1000 ;
	    RECT 57.4000 26.8000 57.8000 27.2000 ;
	    RECT 71.8000 27.1000 72.2000 27.2000 ;
	    RECT 85.4000 27.1000 85.8000 27.2000 ;
	    RECT 89.4000 27.1000 89.8000 27.2000 ;
	    RECT 71.8000 26.8000 89.8000 27.1000 ;
	    RECT 94.2000 27.1000 94.6000 27.2000 ;
	    RECT 107.8000 27.1000 108.2000 27.2000 ;
	    RECT 119.0000 27.1000 119.3000 27.8000 ;
	    RECT 94.2000 26.8000 119.3000 27.1000 ;
	    RECT 127.0000 27.1000 127.4000 27.2000 ;
	    RECT 130.2000 27.1000 130.6000 27.2000 ;
	    RECT 127.0000 26.8000 130.6000 27.1000 ;
	    RECT 7.8000 26.1000 8.2000 26.2000 ;
	    RECT 7.0000 25.8000 8.2000 26.1000 ;
	    RECT 10.2000 26.1000 10.6000 26.2000 ;
	    RECT 17.4000 26.1000 17.8000 26.2000 ;
	    RECT 10.2000 25.8000 17.8000 26.1000 ;
	    RECT 20.6000 25.8000 21.0000 26.2000 ;
	    RECT 31.0000 26.1000 31.3000 26.8000 ;
	    RECT 44.6000 26.1000 45.0000 26.2000 ;
	    RECT 31.0000 25.8000 45.0000 26.1000 ;
	    RECT 50.2000 26.1000 50.6000 26.2000 ;
	    RECT 52.6000 26.1000 53.0000 26.2000 ;
	    RECT 55.0000 26.1000 55.4000 26.2000 ;
	    RECT 50.2000 25.8000 52.1000 26.1000 ;
	    RECT 52.6000 25.8000 55.4000 26.1000 ;
	    RECT 56.6000 26.1000 57.0000 26.2000 ;
	    RECT 57.4000 26.1000 57.7000 26.8000 ;
	    RECT 56.6000 25.8000 57.7000 26.1000 ;
	    RECT 61.4000 25.8000 61.8000 26.2000 ;
	    RECT 63.8000 26.1000 64.2000 26.2000 ;
	    RECT 65.4000 26.1000 65.8000 26.2000 ;
	    RECT 63.8000 25.8000 65.8000 26.1000 ;
	    RECT 75.8000 26.1000 76.2000 26.2000 ;
	    RECT 81.4000 26.1000 81.8000 26.2000 ;
	    RECT 75.8000 25.8000 81.8000 26.1000 ;
	    RECT 82.2000 25.8000 82.6000 26.2000 ;
	    RECT 87.0000 26.1000 87.4000 26.2000 ;
	    RECT 90.2000 26.1000 90.6000 26.2000 ;
	    RECT 103.0000 26.1000 103.4000 26.2000 ;
	    RECT 87.0000 25.8000 103.4000 26.1000 ;
	    RECT 110.2000 26.1000 110.6000 26.2000 ;
	    RECT 115.8000 26.1000 116.2000 26.2000 ;
	    RECT 110.2000 25.8000 116.2000 26.1000 ;
	    RECT 117.4000 26.1000 117.8000 26.2000 ;
	    RECT 127.0000 26.1000 127.4000 26.2000 ;
	    RECT 131.0000 26.1000 131.4000 26.2000 ;
	    RECT 132.6000 26.1000 133.0000 26.2000 ;
	    RECT 117.4000 25.8000 133.0000 26.1000 ;
	    RECT 51.8000 25.2000 52.1000 25.8000 ;
	    RECT 11.8000 25.1000 12.2000 25.2000 ;
	    RECT 12.6000 25.1000 13.0000 25.2000 ;
	    RECT 11.8000 24.8000 13.0000 25.1000 ;
	    RECT 19.0000 25.1000 19.4000 25.2000 ;
	    RECT 39.8000 25.1000 40.2000 25.2000 ;
	    RECT 41.4000 25.1000 41.8000 25.2000 ;
	    RECT 19.0000 24.8000 41.8000 25.1000 ;
	    RECT 51.8000 24.8000 52.2000 25.2000 ;
	    RECT 58.2000 25.1000 58.6000 25.2000 ;
	    RECT 59.8000 25.1000 60.2000 25.2000 ;
	    RECT 58.2000 24.8000 60.2000 25.1000 ;
	    RECT 61.4000 25.1000 61.7000 25.8000 ;
	    RECT 68.6000 25.1000 69.0000 25.2000 ;
	    RECT 61.4000 24.8000 69.0000 25.1000 ;
	    RECT 79.0000 25.1000 79.4000 25.2000 ;
	    RECT 82.2000 25.1000 82.5000 25.8000 ;
	    RECT 83.8000 25.1000 84.2000 25.2000 ;
	    RECT 79.0000 24.8000 84.2000 25.1000 ;
	    RECT 136.6000 25.1000 137.0000 25.2000 ;
	    RECT 145.4000 25.1000 145.8000 25.2000 ;
	    RECT 136.6000 24.8000 145.8000 25.1000 ;
	    RECT 24.6000 24.1000 25.0000 24.2000 ;
	    RECT 32.6000 24.1000 33.0000 24.2000 ;
	    RECT 24.6000 23.8000 33.0000 24.1000 ;
	    RECT 47.8000 24.1000 48.2000 24.2000 ;
	    RECT 49.4000 24.1000 49.8000 24.2000 ;
	    RECT 55.8000 24.1000 56.2000 24.2000 ;
	    RECT 47.8000 23.8000 49.8000 24.1000 ;
	    RECT 55.0000 23.8000 56.2000 24.1000 ;
	    RECT 57.4000 24.1000 57.8000 24.2000 ;
	    RECT 61.4000 24.1000 61.8000 24.2000 ;
	    RECT 57.4000 23.8000 61.8000 24.1000 ;
	    RECT 63.0000 24.1000 63.4000 24.2000 ;
	    RECT 64.6000 24.1000 65.0000 24.2000 ;
	    RECT 63.0000 23.8000 65.0000 24.1000 ;
	    RECT 65.4000 23.8000 65.8000 24.2000 ;
	    RECT 105.4000 24.1000 105.8000 24.2000 ;
	    RECT 114.2000 24.1000 114.6000 24.2000 ;
	    RECT 105.4000 23.8000 114.6000 24.1000 ;
	    RECT 65.4000 23.2000 65.7000 23.8000 ;
	    RECT 31.0000 23.1000 31.4000 23.2000 ;
	    RECT 47.8000 23.1000 48.2000 23.2000 ;
	    RECT 31.0000 22.8000 48.2000 23.1000 ;
	    RECT 48.6000 23.1000 49.0000 23.2000 ;
	    RECT 55.0000 23.1000 55.4000 23.2000 ;
	    RECT 48.6000 22.8000 55.4000 23.1000 ;
	    RECT 65.4000 22.8000 65.8000 23.2000 ;
	    RECT 27.0000 22.1000 27.4000 22.2000 ;
	    RECT 48.6000 22.1000 49.0000 22.2000 ;
	    RECT 27.0000 21.8000 49.0000 22.1000 ;
	    RECT 64.6000 21.2000 64.9000 22.1000 ;
	    RECT 64.6000 20.8000 65.0000 21.2000 ;
	    RECT 65.4000 20.1000 65.8000 20.2000 ;
	    RECT 77.4000 20.1000 77.8000 20.2000 ;
	    RECT 49.4000 19.8000 77.8000 20.1000 ;
	    RECT 11.0000 19.1000 11.4000 19.2000 ;
	    RECT 16.6000 19.1000 17.0000 19.2000 ;
	    RECT 27.8000 19.1000 28.2000 19.2000 ;
	    RECT 11.0000 18.8000 28.2000 19.1000 ;
	    RECT 32.6000 19.1000 33.0000 19.2000 ;
	    RECT 49.4000 19.1000 49.7000 19.8000 ;
	    RECT 32.6000 18.8000 49.7000 19.1000 ;
	    RECT 51.8000 19.1000 52.2000 19.2000 ;
	    RECT 59.0000 19.1000 59.4000 19.2000 ;
	    RECT 51.8000 18.8000 59.4000 19.1000 ;
	    RECT 63.8000 19.1000 64.2000 19.2000 ;
	    RECT 65.4000 19.1000 65.8000 19.2000 ;
	    RECT 63.8000 18.8000 65.8000 19.1000 ;
	    RECT 69.4000 18.8000 69.8000 19.2000 ;
	    RECT 20.6000 18.1000 21.0000 18.2000 ;
	    RECT 28.6000 18.1000 29.0000 18.2000 ;
	    RECT 20.6000 17.8000 29.0000 18.1000 ;
	    RECT 51.8000 18.1000 52.2000 18.2000 ;
	    RECT 52.6000 18.1000 53.0000 18.2000 ;
	    RECT 51.8000 17.8000 53.0000 18.1000 ;
	    RECT 55.0000 18.1000 55.4000 18.2000 ;
	    RECT 69.4000 18.1000 69.7000 18.8000 ;
	    RECT 55.0000 17.8000 69.7000 18.1000 ;
	    RECT 75.0000 18.1000 75.4000 18.2000 ;
	    RECT 94.2000 18.1000 94.6000 18.2000 ;
	    RECT 75.0000 17.8000 94.6000 18.1000 ;
	    RECT 11.0000 17.1000 11.4000 17.2000 ;
	    RECT 13.4000 17.1000 13.8000 17.2000 ;
	    RECT 25.4000 17.1000 25.8000 17.2000 ;
	    RECT 30.2000 17.1000 30.6000 17.2000 ;
	    RECT 11.0000 16.8000 30.6000 17.1000 ;
	    RECT 57.4000 16.8000 57.8000 17.2000 ;
	    RECT 59.0000 17.1000 59.4000 17.2000 ;
	    RECT 60.6000 17.1000 61.0000 17.2000 ;
	    RECT 59.0000 16.8000 61.0000 17.1000 ;
	    RECT 63.0000 17.1000 63.4000 17.2000 ;
	    RECT 83.0000 17.1000 83.4000 17.2000 ;
	    RECT 63.0000 16.8000 83.4000 17.1000 ;
	    RECT 120.6000 17.1000 121.0000 17.2000 ;
	    RECT 143.8000 17.1000 144.2000 17.2000 ;
	    RECT 120.6000 16.8000 144.2000 17.1000 ;
	    RECT 13.4000 15.8000 13.8000 16.2000 ;
	    RECT 16.6000 15.8000 17.0000 16.2000 ;
	    RECT 19.8000 15.8000 20.2000 16.2000 ;
	    RECT 26.2000 16.1000 26.6000 16.2000 ;
	    RECT 31.0000 16.1000 31.4000 16.2000 ;
	    RECT 26.2000 15.8000 31.4000 16.1000 ;
	    RECT 54.2000 16.1000 54.6000 16.2000 ;
	    RECT 57.4000 16.1000 57.7000 16.8000 ;
	    RECT 66.2000 16.1000 66.6000 16.2000 ;
	    RECT 54.2000 15.8000 66.6000 16.1000 ;
	    RECT 87.8000 16.1000 88.2000 16.2000 ;
	    RECT 100.6000 16.1000 101.0000 16.2000 ;
	    RECT 87.8000 15.8000 101.0000 16.1000 ;
	    RECT 110.2000 16.1000 110.6000 16.2000 ;
	    RECT 111.0000 16.1000 111.4000 16.2000 ;
	    RECT 110.2000 15.8000 111.4000 16.1000 ;
	    RECT 121.4000 15.8000 121.8000 16.2000 ;
	    RECT 143.8000 15.8000 144.2000 16.2000 ;
	    RECT 8.6000 15.1000 9.0000 15.2000 ;
	    RECT 13.4000 15.1000 13.7000 15.8000 ;
	    RECT 8.6000 14.8000 13.7000 15.1000 ;
	    RECT 16.6000 15.1000 16.9000 15.8000 ;
	    RECT 19.8000 15.1000 20.1000 15.8000 ;
	    RECT 28.6000 15.2000 28.9000 15.8000 ;
	    RECT 16.6000 14.8000 20.1000 15.1000 ;
	    RECT 22.2000 15.1000 22.6000 15.2000 ;
	    RECT 22.2000 14.8000 24.9000 15.1000 ;
	    RECT 28.6000 14.8000 29.0000 15.2000 ;
	    RECT 35.0000 15.1000 35.4000 15.2000 ;
	    RECT 37.4000 15.1000 37.8000 15.2000 ;
	    RECT 35.0000 14.8000 37.8000 15.1000 ;
	    RECT 39.8000 15.1000 40.2000 15.2000 ;
	    RECT 63.8000 15.1000 64.2000 15.2000 ;
	    RECT 39.8000 14.8000 64.2000 15.1000 ;
	    RECT 64.6000 15.1000 65.0000 15.2000 ;
	    RECT 65.4000 15.1000 65.8000 15.2000 ;
	    RECT 64.6000 14.8000 65.8000 15.1000 ;
	    RECT 71.8000 15.1000 72.2000 15.2000 ;
	    RECT 80.6000 15.1000 81.0000 15.2000 ;
	    RECT 85.4000 15.1000 85.8000 15.2000 ;
	    RECT 71.8000 14.8000 72.9000 15.1000 ;
	    RECT 80.6000 14.8000 85.8000 15.1000 ;
	    RECT 87.0000 15.1000 87.4000 15.2000 ;
	    RECT 101.4000 15.1000 101.8000 15.2000 ;
	    RECT 106.2000 15.1000 106.6000 15.2000 ;
	    RECT 108.6000 15.1000 109.0000 15.2000 ;
	    RECT 110.2000 15.1000 110.6000 15.2000 ;
	    RECT 121.4000 15.1000 121.7000 15.8000 ;
	    RECT 143.8000 15.2000 144.1000 15.8000 ;
	    RECT 87.0000 14.8000 88.1000 15.1000 ;
	    RECT 101.4000 14.8000 121.7000 15.1000 ;
	    RECT 123.0000 15.1000 123.4000 15.2000 ;
	    RECT 128.6000 15.1000 129.0000 15.2000 ;
	    RECT 123.0000 14.8000 129.0000 15.1000 ;
	    RECT 130.2000 15.1000 130.6000 15.2000 ;
	    RECT 130.2000 14.8000 137.7000 15.1000 ;
	    RECT 143.8000 14.8000 144.2000 15.2000 ;
	    RECT 24.6000 14.1000 24.9000 14.8000 ;
	    RECT 137.4000 14.2000 137.7000 14.8000 ;
	    RECT 31.8000 14.1000 32.2000 14.2000 ;
	    RECT 24.6000 13.8000 32.2000 14.1000 ;
	    RECT 68.6000 14.1000 69.0000 14.2000 ;
	    RECT 69.4000 14.1000 69.8000 14.2000 ;
	    RECT 68.6000 13.8000 69.8000 14.1000 ;
	    RECT 71.0000 14.1000 71.4000 14.2000 ;
	    RECT 73.4000 14.1000 73.8000 14.2000 ;
	    RECT 71.0000 13.8000 73.8000 14.1000 ;
	    RECT 81.4000 14.1000 81.8000 14.2000 ;
	    RECT 84.6000 14.1000 85.0000 14.2000 ;
	    RECT 81.4000 13.8000 85.0000 14.1000 ;
	    RECT 89.4000 14.1000 89.8000 14.2000 ;
	    RECT 97.4000 14.1000 97.8000 14.2000 ;
	    RECT 89.4000 13.8000 97.8000 14.1000 ;
	    RECT 137.4000 13.8000 137.8000 14.2000 ;
	    RECT 6.2000 13.1000 6.6000 13.2000 ;
	    RECT 21.4000 13.1000 21.8000 13.2000 ;
	    RECT 6.2000 12.8000 21.8000 13.1000 ;
	    RECT 36.6000 13.1000 37.0000 13.2000 ;
	    RECT 45.4000 13.1000 45.8000 13.2000 ;
	    RECT 36.6000 12.8000 45.8000 13.1000 ;
	    RECT 51.8000 12.8000 52.2000 13.2000 ;
	    RECT 52.6000 13.1000 53.0000 13.2000 ;
	    RECT 59.8000 13.1000 60.2000 13.2000 ;
	    RECT 52.6000 12.8000 60.2000 13.1000 ;
	    RECT 70.2000 13.1000 70.6000 13.2000 ;
	    RECT 78.2000 13.1000 78.6000 13.2000 ;
	    RECT 70.2000 12.8000 78.6000 13.1000 ;
	    RECT 94.2000 13.1000 94.6000 13.2000 ;
	    RECT 95.8000 13.1000 96.2000 13.2000 ;
	    RECT 94.2000 12.8000 96.2000 13.1000 ;
	    RECT 102.2000 12.8000 102.6000 13.2000 ;
	    RECT 110.2000 13.1000 110.6000 13.2000 ;
	    RECT 114.2000 13.1000 114.6000 13.2000 ;
	    RECT 110.2000 12.8000 114.6000 13.1000 ;
	    RECT 51.8000 12.2000 52.1000 12.8000 ;
	    RECT 1.4000 12.1000 1.8000 12.2000 ;
	    RECT 2.2000 12.1000 2.6000 12.2000 ;
	    RECT 1.4000 11.8000 2.6000 12.1000 ;
	    RECT 16.6000 12.1000 17.0000 12.2000 ;
	    RECT 20.6000 12.1000 21.0000 12.2000 ;
	    RECT 16.6000 11.8000 21.0000 12.1000 ;
	    RECT 27.0000 12.1000 27.4000 12.2000 ;
	    RECT 51.0000 12.1000 51.4000 12.2000 ;
	    RECT 27.0000 11.8000 51.4000 12.1000 ;
	    RECT 51.8000 11.8000 52.2000 12.2000 ;
	    RECT 55.0000 12.1000 55.4000 12.2000 ;
	    RECT 55.8000 12.1000 56.2000 12.2000 ;
	    RECT 55.0000 11.8000 56.2000 12.1000 ;
	    RECT 75.0000 12.1000 75.4000 12.2000 ;
	    RECT 86.2000 12.1000 86.6000 12.2000 ;
	    RECT 87.8000 12.1000 88.2000 12.2000 ;
	    RECT 102.2000 12.1000 102.5000 12.8000 ;
	    RECT 75.0000 11.8000 87.3000 12.1000 ;
	    RECT 87.8000 11.8000 102.5000 12.1000 ;
	    RECT 107.0000 11.8000 107.4000 12.2000 ;
	    RECT 131.8000 12.1000 132.2000 12.2000 ;
	    RECT 143.0000 12.1000 143.4000 12.2000 ;
	    RECT 131.8000 11.8000 143.4000 12.1000 ;
	    RECT 107.0000 11.2000 107.3000 11.8000 ;
	    RECT 9.4000 11.1000 9.8000 11.2000 ;
	    RECT 18.2000 11.1000 18.6000 11.2000 ;
	    RECT 9.4000 10.8000 18.6000 11.1000 ;
	    RECT 23.8000 11.1000 24.2000 11.2000 ;
	    RECT 36.6000 11.1000 37.0000 11.2000 ;
	    RECT 39.8000 11.1000 40.2000 11.2000 ;
	    RECT 23.8000 10.8000 40.2000 11.1000 ;
	    RECT 40.6000 11.1000 41.0000 11.2000 ;
	    RECT 43.0000 11.1000 43.4000 11.2000 ;
	    RECT 40.6000 10.8000 43.4000 11.1000 ;
	    RECT 49.4000 11.1000 49.8000 11.2000 ;
	    RECT 51.0000 11.1000 51.4000 11.2000 ;
	    RECT 49.4000 10.8000 51.4000 11.1000 ;
	    RECT 107.0000 10.8000 107.4000 11.2000 ;
	    RECT 18.2000 10.1000 18.6000 10.2000 ;
	    RECT 23.8000 10.1000 24.2000 10.2000 ;
	    RECT 18.2000 9.8000 24.2000 10.1000 ;
	    RECT 35.0000 10.1000 35.4000 10.2000 ;
	    RECT 43.8000 10.1000 44.2000 10.2000 ;
	    RECT 35.0000 9.8000 44.2000 10.1000 ;
	    RECT 83.8000 10.1000 84.2000 10.2000 ;
	    RECT 95.0000 10.1000 95.4000 10.2000 ;
	    RECT 83.8000 9.8000 95.4000 10.1000 ;
	    RECT 7.0000 9.1000 7.4000 9.2000 ;
	    RECT 11.8000 9.1000 12.2000 9.2000 ;
	    RECT 7.0000 8.8000 12.2000 9.1000 ;
	    RECT 15.8000 9.1000 16.2000 9.2000 ;
	    RECT 22.2000 9.1000 22.6000 9.2000 ;
	    RECT 15.8000 8.8000 22.6000 9.1000 ;
	    RECT 29.4000 9.1000 29.8000 9.2000 ;
	    RECT 38.2000 9.1000 38.6000 9.2000 ;
	    RECT 29.4000 8.8000 38.6000 9.1000 ;
	    RECT 41.4000 9.1000 41.8000 9.2000 ;
	    RECT 47.0000 9.1000 47.4000 9.2000 ;
	    RECT 41.4000 8.8000 47.4000 9.1000 ;
	    RECT 53.4000 8.8000 53.8000 9.2000 ;
	    RECT 71.0000 9.1000 71.4000 9.2000 ;
	    RECT 79.8000 9.1000 80.2000 9.2000 ;
	    RECT 103.8000 9.1000 104.2000 9.2000 ;
	    RECT 71.0000 8.8000 80.2000 9.1000 ;
	    RECT 93.4000 8.8000 104.2000 9.1000 ;
	    RECT 8.6000 8.1000 9.0000 8.2000 ;
	    RECT 10.2000 8.1000 10.6000 8.2000 ;
	    RECT 15.8000 8.1000 16.2000 8.2000 ;
	    RECT 8.6000 7.8000 16.2000 8.1000 ;
	    RECT 53.4000 7.8000 53.7000 8.8000 ;
	    RECT 93.4000 8.2000 93.7000 8.8000 ;
	    RECT 55.0000 8.1000 55.4000 8.2000 ;
	    RECT 80.6000 8.1000 81.0000 8.2000 ;
	    RECT 55.0000 7.8000 81.0000 8.1000 ;
	    RECT 81.4000 8.1000 81.8000 8.2000 ;
	    RECT 92.6000 8.1000 93.0000 8.2000 ;
	    RECT 81.4000 7.8000 93.0000 8.1000 ;
	    RECT 93.4000 7.8000 93.8000 8.2000 ;
	    RECT 144.6000 7.8000 145.0000 8.2000 ;
	    RECT 3.8000 7.1000 4.2000 7.2000 ;
	    RECT 11.8000 7.1000 12.2000 7.2000 ;
	    RECT 12.6000 7.1000 13.0000 7.2000 ;
	    RECT 28.6000 7.1000 29.0000 7.2000 ;
	    RECT 29.4000 7.1000 29.8000 7.2000 ;
	    RECT 3.8000 6.8000 8.9000 7.1000 ;
	    RECT 11.8000 6.8000 29.8000 7.1000 ;
	    RECT 43.8000 7.1000 44.2000 7.2000 ;
	    RECT 48.6000 7.1000 49.0000 7.2000 ;
	    RECT 43.8000 6.8000 49.0000 7.1000 ;
	    RECT 51.0000 7.1000 51.4000 7.2000 ;
	    RECT 58.2000 7.1000 58.6000 7.2000 ;
	    RECT 51.0000 6.8000 58.6000 7.1000 ;
	    RECT 69.4000 6.8000 69.8000 7.2000 ;
	    RECT 90.2000 7.1000 90.6000 7.2000 ;
	    RECT 78.2000 6.8000 90.6000 7.1000 ;
	    RECT 107.0000 6.8000 107.4000 7.2000 ;
	    RECT 144.6000 6.8000 144.9000 7.8000 ;
	    RECT 5.4000 6.1000 5.8000 6.2000 ;
	    RECT 7.8000 6.1000 8.2000 6.2000 ;
	    RECT 5.4000 5.8000 8.2000 6.1000 ;
	    RECT 8.6000 6.1000 8.9000 6.8000 ;
	    RECT 18.2000 6.1000 18.6000 6.2000 ;
	    RECT 23.0000 6.1000 23.4000 6.2000 ;
	    RECT 8.6000 5.8000 23.4000 6.1000 ;
	    RECT 29.4000 6.1000 29.8000 6.2000 ;
	    RECT 32.6000 6.1000 33.0000 6.2000 ;
	    RECT 42.2000 6.1000 42.6000 6.2000 ;
	    RECT 53.4000 6.1000 53.8000 6.2000 ;
	    RECT 29.4000 5.8000 42.6000 6.1000 ;
	    RECT 46.2000 5.8000 53.8000 6.1000 ;
	    RECT 62.2000 6.1000 62.6000 6.2000 ;
	    RECT 67.0000 6.1000 67.4000 6.2000 ;
	    RECT 62.2000 5.8000 67.4000 6.1000 ;
	    RECT 69.4000 6.1000 69.7000 6.8000 ;
	    RECT 78.2000 6.2000 78.5000 6.8000 ;
	    RECT 75.0000 6.1000 75.4000 6.2000 ;
	    RECT 69.4000 5.8000 75.4000 6.1000 ;
	    RECT 78.2000 5.8000 78.6000 6.2000 ;
	    RECT 90.2000 6.1000 90.5000 6.8000 ;
	    RECT 103.8000 6.1000 104.2000 6.2000 ;
	    RECT 90.2000 5.8000 104.2000 6.1000 ;
	    RECT 107.0000 6.1000 107.3000 6.8000 ;
	    RECT 108.6000 6.1000 109.0000 6.2000 ;
	    RECT 107.0000 5.8000 109.0000 6.1000 ;
	    RECT 113.4000 6.1000 113.8000 6.2000 ;
	    RECT 115.8000 6.1000 116.2000 6.2000 ;
	    RECT 118.2000 6.1000 118.6000 6.2000 ;
	    RECT 119.8000 6.1000 120.2000 6.2000 ;
	    RECT 121.4000 6.1000 121.8000 6.2000 ;
	    RECT 113.4000 5.8000 121.8000 6.1000 ;
	    RECT 138.2000 6.1000 138.6000 6.2000 ;
	    RECT 140.6000 6.1000 141.0000 6.2000 ;
	    RECT 143.0000 6.1000 143.4000 6.2000 ;
	    RECT 146.2000 6.1000 146.6000 6.2000 ;
	    RECT 138.2000 5.8000 146.6000 6.1000 ;
	    RECT 46.2000 5.2000 46.5000 5.8000 ;
	    RECT 15.8000 5.1000 16.2000 5.2000 ;
	    RECT 19.0000 5.1000 19.4000 5.2000 ;
	    RECT 15.8000 4.8000 19.4000 5.1000 ;
	    RECT 25.4000 5.1000 25.8000 5.2000 ;
	    RECT 43.8000 5.1000 44.2000 5.2000 ;
	    RECT 25.4000 4.8000 44.2000 5.1000 ;
	    RECT 46.2000 4.8000 46.6000 5.2000 ;
	    RECT 51.8000 5.1000 52.2000 5.2000 ;
	    RECT 58.2000 5.1000 58.6000 5.2000 ;
	    RECT 51.0000 4.8000 58.6000 5.1000 ;
	    RECT 63.8000 5.1000 64.2000 5.2000 ;
	    RECT 66.2000 5.1000 66.6000 5.2000 ;
	    RECT 63.8000 4.8000 66.6000 5.1000 ;
	    RECT 31.0000 4.1000 31.4000 4.2000 ;
	    RECT 62.2000 4.1000 62.6000 4.2000 ;
	    RECT 31.0000 3.8000 62.6000 4.1000 ;
	    RECT 69.4000 4.1000 69.8000 4.2000 ;
	    RECT 74.2000 4.1000 74.6000 4.2000 ;
	    RECT 69.4000 3.8000 74.6000 4.1000 ;
	    RECT 96.6000 4.1000 97.0000 4.2000 ;
	    RECT 99.8000 4.1000 100.2000 4.2000 ;
	    RECT 106.2000 4.1000 106.6000 4.2000 ;
	    RECT 96.6000 3.8000 106.6000 4.1000 ;
         LAYER metal4 ;
	    RECT 67.0000 112.8000 67.4000 113.2000 ;
	    RECT 67.0000 105.1000 67.3000 112.8000 ;
	    RECT 88.6000 108.8000 89.0000 109.2000 ;
	    RECT 140.6000 108.8000 141.0000 109.2000 ;
	    RECT 67.8000 105.1000 68.2000 105.2000 ;
	    RECT 67.0000 104.8000 68.2000 105.1000 ;
	    RECT 15.0000 89.8000 15.4000 90.2000 ;
	    RECT 72.6000 90.1000 73.0000 90.2000 ;
	    RECT 71.8000 89.8000 73.0000 90.1000 ;
	    RECT 15.0000 47.2000 15.3000 89.8000 ;
	    RECT 17.4000 87.1000 17.8000 87.2000 ;
	    RECT 17.4000 86.8000 18.5000 87.1000 ;
	    RECT 18.2000 74.2000 18.5000 86.8000 ;
	    RECT 71.0000 80.8000 71.4000 81.2000 ;
	    RECT 70.2000 78.8000 70.6000 79.2000 ;
	    RECT 30.2000 75.1000 30.6000 75.2000 ;
	    RECT 29.4000 74.8000 30.6000 75.1000 ;
	    RECT 18.2000 73.8000 18.6000 74.2000 ;
	    RECT 29.4000 58.2000 29.7000 74.8000 ;
	    RECT 70.2000 68.2000 70.5000 78.8000 ;
	    RECT 70.2000 67.8000 70.6000 68.2000 ;
	    RECT 43.0000 66.8000 43.4000 67.2000 ;
	    RECT 29.4000 57.8000 29.8000 58.2000 ;
	    RECT 43.0000 54.2000 43.3000 66.8000 ;
	    RECT 71.0000 66.2000 71.3000 80.8000 ;
	    RECT 71.0000 65.8000 71.4000 66.2000 ;
	    RECT 71.8000 61.2000 72.1000 89.8000 ;
	    RECT 87.0000 89.1000 87.4000 89.2000 ;
	    RECT 87.0000 88.8000 88.1000 89.1000 ;
	    RECT 87.8000 86.2000 88.1000 88.8000 ;
	    RECT 87.8000 85.8000 88.2000 86.2000 ;
	    RECT 72.6000 80.8000 73.0000 81.2000 ;
	    RECT 72.6000 62.2000 72.9000 80.8000 ;
	    RECT 88.6000 67.1000 88.9000 108.8000 ;
	    RECT 139.0000 108.1000 139.4000 108.2000 ;
	    RECT 138.2000 107.8000 139.4000 108.1000 ;
	    RECT 135.0000 105.8000 135.4000 106.2000 ;
	    RECT 120.6000 105.1000 121.0000 105.2000 ;
	    RECT 120.6000 104.8000 121.7000 105.1000 ;
	    RECT 112.6000 89.8000 113.0000 90.2000 ;
	    RECT 93.4000 87.8000 93.8000 88.2000 ;
	    RECT 90.2000 68.8000 90.6000 69.2000 ;
	    RECT 90.2000 67.2000 90.5000 68.8000 ;
	    RECT 89.4000 67.1000 89.8000 67.2000 ;
	    RECT 88.6000 66.8000 89.8000 67.1000 ;
	    RECT 90.2000 66.8000 90.6000 67.2000 ;
	    RECT 72.6000 61.8000 73.0000 62.2000 ;
	    RECT 71.8000 60.8000 72.2000 61.2000 ;
	    RECT 91.0000 56.1000 91.4000 56.2000 ;
	    RECT 90.2000 55.8000 91.4000 56.1000 ;
	    RECT 43.0000 53.8000 43.4000 54.2000 ;
	    RECT 89.4000 52.8000 89.8000 53.2000 ;
	    RECT 89.4000 52.2000 89.7000 52.8000 ;
	    RECT 89.4000 51.8000 89.8000 52.2000 ;
	    RECT 89.4000 49.8000 89.8000 50.2000 ;
	    RECT 15.0000 46.8000 15.4000 47.2000 ;
	    RECT 75.0000 46.8000 75.4000 47.2000 ;
	    RECT 29.4000 43.8000 29.8000 44.2000 ;
	    RECT 27.0000 35.1000 27.4000 35.2000 ;
	    RECT 28.6000 35.1000 29.0000 35.2000 ;
	    RECT 27.0000 34.8000 29.0000 35.1000 ;
	    RECT 19.8000 27.1000 20.2000 27.2000 ;
	    RECT 19.8000 26.8000 20.9000 27.1000 ;
	    RECT 7.8000 26.1000 8.2000 26.2000 ;
	    RECT 7.0000 25.8000 8.2000 26.1000 ;
	    RECT 12.6000 25.1000 13.0000 25.2000 ;
	    RECT 11.8000 24.8000 13.0000 25.1000 ;
	    RECT 11.8000 7.2000 12.1000 24.8000 ;
	    RECT 20.6000 12.2000 20.9000 26.8000 ;
	    RECT 20.6000 11.8000 21.0000 12.2000 ;
	    RECT 29.4000 7.2000 29.7000 43.8000 ;
	    RECT 47.0000 35.1000 47.4000 35.2000 ;
	    RECT 47.8000 35.1000 48.2000 35.2000 ;
	    RECT 47.0000 34.8000 48.2000 35.1000 ;
	    RECT 53.4000 30.8000 53.8000 31.2000 ;
	    RECT 51.8000 27.8000 52.2000 28.2000 ;
	    RECT 45.4000 26.8000 45.8000 27.2000 ;
	    RECT 45.4000 26.2000 45.7000 26.8000 ;
	    RECT 45.4000 25.8000 45.8000 26.2000 ;
	    RECT 41.4000 24.8000 41.8000 25.2000 ;
	    RECT 39.8000 14.8000 40.2000 15.2000 ;
	    RECT 39.8000 11.2000 40.1000 14.8000 ;
	    RECT 39.8000 10.8000 40.2000 11.2000 ;
	    RECT 41.4000 9.2000 41.7000 24.8000 ;
	    RECT 51.8000 18.2000 52.1000 27.8000 ;
	    RECT 51.8000 17.8000 52.2000 18.2000 ;
	    RECT 51.8000 14.8000 52.2000 15.2000 ;
	    RECT 51.8000 13.2000 52.1000 14.8000 ;
	    RECT 51.8000 12.8000 52.2000 13.2000 ;
	    RECT 51.0000 11.8000 51.4000 12.2000 ;
	    RECT 41.4000 8.8000 41.8000 9.2000 ;
	    RECT 51.0000 7.2000 51.3000 11.8000 ;
	    RECT 53.4000 9.2000 53.7000 30.8000 ;
	    RECT 63.8000 28.8000 64.2000 29.2000 ;
	    RECT 55.0000 26.1000 55.4000 26.2000 ;
	    RECT 55.8000 26.1000 56.2000 26.2000 ;
	    RECT 55.0000 25.8000 56.2000 26.1000 ;
	    RECT 55.8000 24.1000 56.2000 24.2000 ;
	    RECT 55.0000 23.8000 56.2000 24.1000 ;
	    RECT 63.8000 24.1000 64.1000 28.8000 ;
	    RECT 65.4000 26.1000 65.8000 26.2000 ;
	    RECT 64.6000 25.8000 65.8000 26.1000 ;
	    RECT 64.6000 25.2000 64.9000 25.8000 ;
	    RECT 64.6000 24.8000 65.0000 25.2000 ;
	    RECT 64.6000 24.1000 65.0000 24.2000 ;
	    RECT 63.8000 23.8000 65.0000 24.1000 ;
	    RECT 55.0000 12.2000 55.3000 23.8000 ;
	    RECT 65.4000 22.8000 65.8000 23.2000 ;
	    RECT 64.6000 20.8000 65.0000 21.2000 ;
	    RECT 64.6000 15.2000 64.9000 20.8000 ;
	    RECT 65.4000 19.2000 65.7000 22.8000 ;
	    RECT 65.4000 18.8000 65.8000 19.2000 ;
	    RECT 75.0000 18.2000 75.3000 46.8000 ;
	    RECT 89.4000 36.2000 89.7000 49.8000 ;
	    RECT 89.4000 35.8000 89.8000 36.2000 ;
	    RECT 90.2000 26.2000 90.5000 55.8000 ;
	    RECT 91.8000 53.1000 92.2000 53.2000 ;
	    RECT 92.6000 53.1000 93.0000 53.2000 ;
	    RECT 91.8000 52.8000 93.0000 53.1000 ;
	    RECT 91.0000 48.8000 91.4000 49.2000 ;
	    RECT 93.4000 49.1000 93.7000 87.8000 ;
	    RECT 112.6000 80.2000 112.9000 89.8000 ;
	    RECT 119.0000 85.8000 119.4000 86.2000 ;
	    RECT 112.6000 79.8000 113.0000 80.2000 ;
	    RECT 112.6000 78.1000 113.0000 78.2000 ;
	    RECT 113.4000 78.1000 113.8000 78.2000 ;
	    RECT 112.6000 77.8000 113.8000 78.1000 ;
	    RECT 114.2000 78.1000 114.6000 78.2000 ;
	    RECT 115.0000 78.1000 115.4000 78.2000 ;
	    RECT 114.2000 77.8000 115.4000 78.1000 ;
	    RECT 97.4000 76.8000 97.8000 77.2000 ;
	    RECT 97.4000 72.2000 97.7000 76.8000 ;
	    RECT 115.8000 75.8000 116.2000 76.2000 ;
	    RECT 115.8000 73.2000 116.1000 75.8000 ;
	    RECT 115.8000 72.8000 116.2000 73.2000 ;
	    RECT 96.6000 71.8000 97.0000 72.2000 ;
	    RECT 97.4000 71.8000 97.8000 72.2000 ;
	    RECT 96.6000 65.2000 96.9000 71.8000 ;
	    RECT 109.4000 69.8000 109.8000 70.2000 ;
	    RECT 96.6000 64.8000 97.0000 65.2000 ;
	    RECT 109.4000 65.1000 109.7000 69.8000 ;
	    RECT 110.2000 65.1000 110.6000 65.2000 ;
	    RECT 109.4000 64.8000 110.6000 65.1000 ;
	    RECT 118.2000 65.1000 118.6000 65.2000 ;
	    RECT 119.0000 65.1000 119.3000 85.8000 ;
	    RECT 118.2000 64.8000 119.3000 65.1000 ;
	    RECT 101.4000 56.1000 101.8000 56.2000 ;
	    RECT 102.2000 56.1000 102.6000 56.2000 ;
	    RECT 101.4000 55.8000 102.6000 56.1000 ;
	    RECT 94.2000 49.1000 94.6000 49.2000 ;
	    RECT 93.4000 48.8000 94.6000 49.1000 ;
	    RECT 91.0000 47.2000 91.3000 48.8000 ;
	    RECT 91.0000 46.8000 91.4000 47.2000 ;
	    RECT 91.8000 44.8000 92.2000 45.2000 ;
	    RECT 95.0000 45.1000 95.4000 45.2000 ;
	    RECT 95.0000 44.8000 96.1000 45.1000 ;
	    RECT 91.8000 44.2000 92.1000 44.8000 ;
	    RECT 91.8000 43.8000 92.2000 44.2000 ;
	    RECT 103.0000 40.8000 103.4000 41.2000 ;
	    RECT 103.0000 26.2000 103.3000 40.8000 ;
	    RECT 107.0000 33.8000 107.4000 34.2000 ;
	    RECT 90.2000 25.8000 90.6000 26.2000 ;
	    RECT 103.0000 25.8000 103.4000 26.2000 ;
	    RECT 75.0000 17.8000 75.4000 18.2000 ;
	    RECT 64.6000 14.8000 65.0000 15.2000 ;
	    RECT 71.8000 15.1000 72.2000 15.2000 ;
	    RECT 87.0000 15.1000 87.4000 15.2000 ;
	    RECT 71.8000 14.8000 72.9000 15.1000 ;
	    RECT 87.0000 14.8000 88.1000 15.1000 ;
	    RECT 87.8000 14.2000 88.1000 14.8000 ;
	    RECT 69.4000 14.1000 69.8000 14.2000 ;
	    RECT 70.2000 14.1000 70.6000 14.2000 ;
	    RECT 69.4000 13.8000 70.6000 14.1000 ;
	    RECT 87.8000 13.8000 88.2000 14.2000 ;
	    RECT 107.0000 12.2000 107.3000 33.8000 ;
	    RECT 110.2000 16.2000 110.5000 64.8000 ;
	    RECT 121.4000 61.2000 121.7000 104.8000 ;
	    RECT 135.0000 72.2000 135.3000 105.8000 ;
	    RECT 137.4000 76.1000 137.8000 76.2000 ;
	    RECT 136.6000 75.8000 137.8000 76.1000 ;
	    RECT 127.0000 71.8000 127.4000 72.2000 ;
	    RECT 135.0000 71.8000 135.4000 72.2000 ;
	    RECT 127.0000 66.2000 127.3000 71.8000 ;
	    RECT 127.8000 70.8000 128.2000 71.2000 ;
	    RECT 127.0000 65.8000 127.4000 66.2000 ;
	    RECT 127.8000 66.1000 128.1000 70.8000 ;
	    RECT 128.6000 66.1000 129.0000 66.2000 ;
	    RECT 127.8000 65.8000 129.0000 66.1000 ;
	    RECT 121.4000 60.8000 121.8000 61.2000 ;
	    RECT 123.8000 58.1000 124.2000 58.2000 ;
	    RECT 123.8000 57.8000 124.9000 58.1000 ;
	    RECT 113.4000 56.1000 113.8000 56.2000 ;
	    RECT 113.4000 55.8000 114.5000 56.1000 ;
	    RECT 124.6000 53.2000 124.9000 57.8000 ;
	    RECT 124.6000 52.8000 125.0000 53.2000 ;
	    RECT 127.0000 27.2000 127.3000 65.8000 ;
	    RECT 127.0000 26.8000 127.4000 27.2000 ;
	    RECT 136.6000 25.2000 136.9000 75.8000 ;
	    RECT 138.2000 44.2000 138.5000 107.8000 ;
	    RECT 138.2000 43.8000 138.6000 44.2000 ;
	    RECT 140.6000 35.2000 140.9000 108.8000 ;
	    RECT 143.8000 80.8000 144.2000 81.2000 ;
	    RECT 140.6000 34.8000 141.0000 35.2000 ;
	    RECT 136.6000 24.8000 137.0000 25.2000 ;
	    RECT 143.8000 17.2000 144.1000 80.8000 ;
	    RECT 144.6000 54.8000 145.0000 55.2000 ;
	    RECT 143.8000 16.8000 144.2000 17.2000 ;
	    RECT 143.8000 16.2000 144.1000 16.8000 ;
	    RECT 110.2000 15.8000 110.6000 16.2000 ;
	    RECT 143.8000 15.8000 144.2000 16.2000 ;
	    RECT 55.0000 11.8000 55.4000 12.2000 ;
	    RECT 107.0000 11.8000 107.4000 12.2000 ;
	    RECT 53.4000 8.8000 53.8000 9.2000 ;
	    RECT 144.6000 8.2000 144.9000 54.8000 ;
	    RECT 144.6000 7.8000 145.0000 8.2000 ;
	    RECT 11.8000 6.8000 12.2000 7.2000 ;
	    RECT 29.4000 6.8000 29.8000 7.2000 ;
	    RECT 51.0000 6.8000 51.4000 7.2000 ;
         LAYER metal5 ;
	    RECT 113.4000 78.1000 113.8000 78.2000 ;
	    RECT 114.2000 78.1000 114.6000 78.2000 ;
	    RECT 113.4000 77.8000 114.6000 78.1000 ;
	    RECT 102.2000 56.1000 102.6000 56.2000 ;
	    RECT 113.4000 56.1000 113.8000 56.2000 ;
	    RECT 102.2000 55.8000 113.8000 56.1000 ;
	    RECT 89.4000 53.1000 89.8000 53.2000 ;
	    RECT 91.8000 53.1000 92.2000 53.2000 ;
	    RECT 89.4000 52.8000 92.2000 53.1000 ;
	    RECT 91.8000 45.1000 92.2000 45.2000 ;
	    RECT 95.0000 45.1000 95.4000 45.2000 ;
	    RECT 91.8000 44.8000 95.4000 45.1000 ;
	    RECT 28.6000 35.1000 29.0000 35.2000 ;
	    RECT 47.0000 35.1000 47.4000 35.2000 ;
	    RECT 28.6000 34.8000 47.4000 35.1000 ;
	    RECT 7.8000 26.1000 8.2000 26.2000 ;
	    RECT 45.4000 26.1000 45.8000 26.2000 ;
	    RECT 7.8000 25.8000 45.8000 26.1000 ;
	    RECT 55.8000 26.1000 56.2000 26.2000 ;
	    RECT 55.8000 25.8000 64.9000 26.1000 ;
	    RECT 64.6000 25.2000 64.9000 25.8000 ;
	    RECT 64.6000 24.8000 65.0000 25.2000 ;
	    RECT 51.8000 15.1000 52.2000 15.2000 ;
	    RECT 71.8000 15.1000 72.2000 15.2000 ;
	    RECT 51.8000 14.8000 72.2000 15.1000 ;
	    RECT 70.2000 14.1000 70.6000 14.2000 ;
	    RECT 87.8000 14.1000 88.2000 14.2000 ;
	    RECT 70.2000 13.8000 88.2000 14.1000 ;
   END
END BFCPU
