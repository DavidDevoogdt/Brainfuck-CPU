magic
tech scmos
timestamp 1537603335
<< metal1 >>
rect 476 1203 477 1207
rect 481 1203 482 1207
rect 486 1203 488 1207
rect 478 1188 494 1191
rect 1086 1168 1094 1171
rect 1470 1168 1486 1171
rect 662 1161 665 1168
rect 1086 1166 1090 1168
rect 1110 1166 1114 1168
rect 662 1158 673 1161
rect 118 1148 129 1151
rect 126 1142 129 1148
rect 390 1148 398 1151
rect 430 1148 441 1151
rect 538 1148 569 1151
rect 620 1148 638 1151
rect 798 1151 802 1153
rect 438 1142 441 1148
rect 798 1148 809 1151
rect 998 1148 1022 1151
rect 1206 1151 1210 1153
rect 1262 1151 1266 1153
rect 1170 1148 1177 1151
rect 1206 1148 1217 1151
rect 1254 1148 1266 1151
rect 574 1138 593 1141
rect 638 1138 646 1141
rect 998 1138 1001 1148
rect 1398 1148 1406 1151
rect 782 1133 786 1138
rect 442 1128 449 1131
rect 1278 1131 1282 1136
rect 1278 1128 1294 1131
rect 338 1118 340 1122
rect 980 1118 982 1122
rect 980 1103 981 1107
rect 985 1103 986 1107
rect 990 1103 992 1107
rect 562 1088 569 1091
rect 46 1078 62 1081
rect 134 1078 145 1081
rect 46 1074 50 1078
rect 206 1072 210 1077
rect 406 1071 409 1081
rect 386 1068 409 1071
rect 446 1068 457 1071
rect 478 1068 502 1071
rect 540 1068 550 1071
rect 22 1058 34 1061
rect 62 1058 70 1061
rect 142 1061 145 1068
rect 142 1058 153 1061
rect 182 1058 194 1061
rect 222 1058 230 1061
rect 290 1058 305 1061
rect 374 1058 406 1061
rect 506 1058 529 1061
rect 614 1058 622 1061
rect 646 1061 649 1071
rect 674 1068 681 1071
rect 726 1068 737 1071
rect 926 1068 929 1078
rect 1246 1071 1249 1081
rect 1218 1068 1233 1071
rect 1246 1068 1265 1071
rect 1334 1071 1337 1081
rect 1334 1068 1353 1071
rect 646 1058 665 1061
rect 708 1058 726 1061
rect 1126 1058 1153 1061
rect 1362 1058 1369 1061
rect 1374 1058 1382 1061
rect 30 1057 34 1058
rect 190 1057 194 1058
rect 562 1048 569 1051
rect 658 1038 665 1041
rect 746 1038 753 1041
rect 1290 1038 1291 1042
rect 1114 1018 1115 1022
rect 1194 1018 1195 1022
rect 476 1003 477 1007
rect 481 1003 482 1007
rect 486 1003 488 1007
rect 450 988 451 992
rect 893 988 894 992
rect 954 988 955 992
rect 1462 988 1486 991
rect 74 968 77 972
rect 1258 968 1259 972
rect 462 958 489 961
rect 1162 958 1166 962
rect 54 951 58 953
rect 46 948 58 951
rect 338 948 345 951
rect 410 948 414 951
rect 670 948 678 951
rect 706 948 713 951
rect 1022 951 1026 953
rect 958 948 969 951
rect 1014 948 1026 951
rect 1166 948 1174 951
rect 1206 948 1217 951
rect 93 938 94 942
rect 62 936 66 938
rect 182 932 185 942
rect 422 938 441 941
rect 1178 938 1185 941
rect 1214 938 1217 948
rect 1378 938 1385 941
rect 574 931 577 938
rect 1038 932 1042 936
rect 574 928 585 931
rect 646 928 657 931
rect 694 928 705 931
rect 378 918 380 922
rect 980 903 981 907
rect 985 903 986 907
rect 990 903 992 907
rect 146 888 148 892
rect 586 888 588 892
rect 756 888 758 892
rect 46 874 50 878
rect 482 868 489 871
rect 562 868 566 871
rect 686 868 697 871
rect 894 868 905 871
rect 950 868 958 871
rect 1042 868 1049 871
rect 1318 868 1330 871
rect 1470 868 1486 871
rect 22 858 34 861
rect 694 862 697 868
rect 254 858 265 861
rect 506 858 510 861
rect 546 858 553 861
rect 658 858 673 861
rect 902 861 905 868
rect 902 858 913 861
rect 1054 858 1078 861
rect 1134 861 1138 864
rect 1126 858 1138 861
rect 30 857 34 858
rect 482 848 489 851
rect 642 848 649 851
rect 306 838 308 842
rect 802 838 805 842
rect 194 818 195 822
rect 476 803 477 807
rect 481 803 482 807
rect 486 803 488 807
rect 437 788 438 792
rect 740 788 742 792
rect 1306 788 1307 792
rect 1454 788 1486 791
rect 1086 772 1089 781
rect 118 768 129 771
rect 126 762 129 768
rect 190 768 217 771
rect 1146 768 1147 772
rect 1386 768 1387 772
rect 158 761 161 768
rect 150 758 161 761
rect 474 758 494 761
rect 994 758 1017 761
rect 1398 758 1409 761
rect 22 748 38 751
rect 66 748 89 751
rect 318 748 337 751
rect 342 748 353 751
rect 582 751 586 752
rect 566 748 586 751
rect 86 741 89 748
rect 86 738 94 741
rect 566 742 569 748
rect 1094 751 1098 754
rect 1094 748 1113 751
rect 1234 748 1241 751
rect 1286 748 1297 751
rect 410 738 417 741
rect 422 738 430 741
rect 502 738 510 741
rect 758 738 777 741
rect 1050 738 1062 741
rect 1294 738 1297 748
rect 1366 738 1377 741
rect 66 728 73 731
rect 534 728 542 731
rect 470 718 478 721
rect 802 718 803 722
rect 980 703 981 707
rect 985 703 986 707
rect 990 703 992 707
rect 969 688 998 691
rect 1006 688 1017 691
rect 1142 688 1150 691
rect 1470 688 1486 691
rect 1006 682 1009 688
rect 222 678 233 681
rect 898 678 910 681
rect 46 672 50 677
rect 134 668 145 671
rect 562 668 569 671
rect 590 668 601 671
rect 606 668 614 671
rect 782 668 806 671
rect 930 668 953 671
rect 1038 668 1046 671
rect 1410 668 1417 671
rect 22 658 34 661
rect 142 662 145 668
rect 378 658 393 661
rect 478 658 486 661
rect 554 658 566 661
rect 570 658 577 661
rect 706 658 713 661
rect 914 658 921 661
rect 1050 658 1057 661
rect 1254 658 1262 661
rect 1350 658 1358 661
rect 30 657 34 658
rect 370 648 374 652
rect 446 648 457 651
rect 1042 648 1049 651
rect 1414 651 1417 658
rect 1414 648 1425 651
rect 278 638 298 641
rect 1066 638 1073 641
rect 1182 638 1209 641
rect 278 628 281 638
rect 309 618 310 622
rect 476 603 477 607
rect 481 603 482 607
rect 486 603 488 607
rect 1194 588 1195 592
rect 114 568 117 572
rect 1133 568 1134 572
rect 1258 568 1259 572
rect 1294 566 1298 568
rect 1422 566 1426 568
rect 1470 568 1478 571
rect 1470 566 1474 568
rect 638 558 657 561
rect 214 548 222 551
rect 546 548 553 551
rect 754 548 761 551
rect 838 551 841 561
rect 818 548 825 551
rect 838 548 857 551
rect 878 548 889 551
rect 1174 548 1185 551
rect 1206 551 1209 561
rect 1270 558 1289 561
rect 1206 548 1225 551
rect 1230 548 1238 551
rect 1378 548 1385 551
rect 1426 548 1433 551
rect 370 538 377 541
rect 606 538 625 541
rect 638 538 646 541
rect 682 538 689 541
rect 742 538 750 541
rect 786 538 793 541
rect 862 538 870 541
rect 1146 538 1153 541
rect 1182 538 1185 548
rect 1350 538 1369 541
rect 722 528 737 531
rect 762 528 769 531
rect 1330 528 1337 531
rect 514 518 516 522
rect 1418 518 1419 522
rect 980 503 981 507
rect 985 503 986 507
rect 990 503 992 507
rect 706 478 713 482
rect 742 478 750 481
rect 982 478 1017 481
rect 550 474 554 478
rect 710 472 713 478
rect 102 468 113 471
rect 178 468 185 471
rect 454 468 482 471
rect 642 468 649 471
rect 654 468 670 471
rect 766 468 785 471
rect 966 468 977 471
rect 1294 471 1297 481
rect 1462 478 1470 481
rect 1294 468 1313 471
rect 1366 468 1377 471
rect 102 462 105 468
rect 254 461 257 468
rect 238 458 257 461
rect 966 462 969 468
rect 1206 458 1214 461
rect 294 448 302 451
rect 334 448 342 451
rect 630 448 641 451
rect 710 448 721 451
rect 798 448 806 451
rect 854 448 873 451
rect 258 438 265 441
rect 326 438 353 441
rect 885 438 886 442
rect 957 438 958 442
rect 1050 438 1053 442
rect 1341 418 1342 422
rect 476 403 477 407
rect 481 403 482 407
rect 486 403 488 407
rect 1454 368 1486 371
rect 470 358 497 361
rect 1046 358 1054 361
rect 30 351 34 353
rect 22 348 34 351
rect 142 348 153 351
rect 298 348 310 351
rect 462 351 465 358
rect 378 348 385 351
rect 462 348 473 351
rect 514 348 518 351
rect 530 348 537 351
rect 542 348 569 351
rect 618 348 625 351
rect 850 348 865 351
rect 966 348 982 351
rect 1078 348 1089 351
rect 142 342 145 348
rect 294 338 321 341
rect 646 338 681 341
rect 790 338 809 341
rect 822 338 841 341
rect 870 338 889 341
rect 910 338 918 341
rect 946 338 953 341
rect 994 338 1001 341
rect 1086 338 1089 348
rect 46 331 50 336
rect 46 328 62 331
rect 134 328 145 331
rect 294 328 297 338
rect 338 328 345 331
rect 350 328 361 331
rect 710 328 734 331
rect 772 328 785 331
rect 822 328 825 338
rect 918 328 929 331
rect 1366 328 1385 331
rect 710 322 713 328
rect 178 318 179 322
rect 450 318 451 322
rect 654 318 662 321
rect 980 303 981 307
rect 985 303 986 307
rect 990 303 992 307
rect 974 288 982 291
rect 326 278 353 281
rect 666 278 673 281
rect 838 278 854 281
rect 1150 278 1161 281
rect 1326 278 1345 281
rect 126 268 145 271
rect 150 268 166 271
rect 198 268 206 271
rect 370 268 377 271
rect 382 268 390 271
rect 430 268 438 271
rect 510 268 518 271
rect 538 268 548 271
rect 722 268 729 271
rect 1470 268 1486 271
rect 190 258 198 261
rect 322 258 345 261
rect 430 261 434 264
rect 430 258 441 261
rect 446 258 454 261
rect 502 258 510 261
rect 526 258 534 261
rect 578 258 585 261
rect 730 258 737 261
rect 770 258 777 261
rect 986 258 1001 261
rect 1158 261 1161 268
rect 1158 258 1169 261
rect 1214 258 1230 261
rect 498 248 502 252
rect 734 248 745 251
rect 754 248 758 252
rect 570 238 578 241
rect 117 218 118 222
rect 476 203 477 207
rect 481 203 482 207
rect 486 203 488 207
rect 549 188 550 192
rect 426 168 430 171
rect 434 168 441 171
rect 1250 168 1257 171
rect 242 158 249 161
rect 394 158 401 161
rect 418 158 425 161
rect 694 158 705 161
rect 342 148 358 151
rect 374 148 385 151
rect 462 148 505 151
rect 550 148 558 151
rect 574 148 585 151
rect 606 148 617 151
rect 730 148 753 151
rect 778 148 814 151
rect 914 148 921 151
rect 1142 148 1150 151
rect 1222 148 1233 151
rect 1298 148 1313 151
rect 318 141 321 148
rect 374 142 377 148
rect 318 138 329 141
rect 686 141 689 148
rect 1230 142 1233 148
rect 670 138 689 141
rect 850 138 873 141
rect 1030 138 1049 141
rect 1090 138 1097 141
rect 1106 138 1129 141
rect 1166 138 1174 141
rect 1342 138 1354 141
rect 454 131 457 138
rect 394 128 406 131
rect 454 128 465 131
rect 682 128 689 131
rect 742 128 750 131
rect 794 128 801 131
rect 858 128 865 131
rect 958 131 961 138
rect 958 128 974 131
rect 1030 128 1033 138
rect 1070 128 1089 131
rect 1230 128 1241 131
rect 980 103 981 107
rect 985 103 986 107
rect 990 103 992 107
rect 249 88 270 91
rect 434 88 441 91
rect 1300 88 1302 92
rect 1458 88 1459 92
rect 102 78 110 82
rect 102 72 105 78
rect 38 68 46 71
rect 166 68 182 71
rect 358 68 377 71
rect 538 68 545 71
rect 78 61 81 68
rect 38 58 49 61
rect 78 58 89 61
rect 286 58 302 61
rect 358 61 361 68
rect 318 58 337 61
rect 342 58 361 61
rect 446 58 457 61
rect 474 58 505 61
rect 518 58 526 61
rect 622 61 625 68
rect 586 58 601 61
rect 606 58 625 61
rect 934 58 945 61
rect 1038 58 1046 61
rect 1318 61 1321 68
rect 1318 58 1329 61
rect 1366 58 1374 61
rect 318 48 321 58
rect 518 48 521 58
rect 638 51 641 58
rect 934 57 938 58
rect 630 48 641 51
rect 1462 48 1486 51
rect 476 3 477 7
rect 481 3 482 7
rect 486 3 488 7
<< m2contact >>
rect 472 1203 476 1207
rect 477 1203 481 1207
rect 482 1203 486 1207
rect 102 1188 106 1192
rect 214 1188 218 1192
rect 494 1188 498 1192
rect 702 1188 706 1192
rect 822 1188 826 1192
rect 846 1188 850 1192
rect 870 1188 874 1192
rect 894 1188 898 1192
rect 918 1188 922 1192
rect 942 1188 946 1192
rect 1038 1188 1042 1192
rect 1062 1188 1066 1192
rect 1230 1188 1234 1192
rect 1238 1188 1242 1192
rect 1374 1188 1378 1192
rect 1422 1188 1426 1192
rect 1446 1188 1450 1192
rect 6 1168 10 1172
rect 222 1168 226 1172
rect 662 1168 666 1172
rect 1094 1168 1098 1172
rect 1110 1168 1114 1172
rect 1486 1168 1490 1172
rect 398 1158 402 1162
rect 646 1158 650 1162
rect 70 1147 74 1151
rect 142 1148 146 1152
rect 198 1148 202 1152
rect 254 1148 258 1152
rect 286 1147 290 1151
rect 382 1148 386 1152
rect 398 1148 402 1152
rect 406 1148 410 1152
rect 462 1148 466 1152
rect 534 1148 538 1152
rect 638 1148 642 1152
rect 686 1148 690 1152
rect 734 1147 738 1151
rect 830 1148 834 1152
rect 854 1148 858 1152
rect 878 1148 882 1152
rect 902 1148 906 1152
rect 926 1148 930 1152
rect 1022 1148 1026 1152
rect 1046 1148 1050 1152
rect 1150 1148 1154 1152
rect 1166 1148 1170 1152
rect 1294 1148 1298 1152
rect 126 1138 130 1142
rect 174 1138 178 1142
rect 318 1138 322 1142
rect 366 1138 370 1142
rect 374 1138 378 1142
rect 414 1138 418 1142
rect 438 1138 442 1142
rect 542 1138 546 1142
rect 646 1138 650 1142
rect 662 1138 666 1142
rect 678 1138 682 1142
rect 750 1138 754 1142
rect 782 1138 786 1142
rect 950 1138 954 1142
rect 1326 1147 1330 1151
rect 1358 1148 1362 1152
rect 1406 1148 1410 1152
rect 1430 1148 1434 1152
rect 1454 1148 1458 1152
rect 1070 1138 1074 1142
rect 1094 1138 1098 1142
rect 1126 1138 1130 1142
rect 70 1128 74 1132
rect 182 1128 186 1132
rect 430 1128 434 1132
rect 438 1128 442 1132
rect 454 1128 458 1132
rect 550 1128 554 1132
rect 582 1128 586 1132
rect 1294 1128 1298 1132
rect 190 1118 194 1122
rect 334 1118 338 1122
rect 526 1118 530 1122
rect 646 1118 650 1122
rect 982 1118 986 1122
rect 1086 1118 1090 1122
rect 1110 1118 1114 1122
rect 1206 1118 1210 1122
rect 976 1103 980 1107
rect 981 1103 985 1107
rect 986 1103 990 1107
rect 166 1088 170 1092
rect 382 1088 386 1092
rect 422 1088 426 1092
rect 558 1088 562 1092
rect 598 1088 602 1092
rect 630 1088 634 1092
rect 862 1088 866 1092
rect 958 1088 962 1092
rect 1070 1088 1074 1092
rect 1238 1088 1242 1092
rect 1326 1088 1330 1092
rect 1478 1088 1482 1092
rect 62 1078 66 1082
rect 126 1078 130 1082
rect 254 1078 258 1082
rect 390 1078 394 1082
rect 6 1068 10 1072
rect 142 1068 146 1072
rect 206 1068 210 1072
rect 286 1068 290 1072
rect 334 1068 338 1072
rect 382 1068 386 1072
rect 510 1078 514 1082
rect 742 1078 746 1082
rect 926 1078 930 1082
rect 1078 1078 1082 1082
rect 1086 1078 1090 1082
rect 414 1068 418 1072
rect 502 1068 506 1072
rect 518 1068 522 1072
rect 550 1068 554 1072
rect 590 1068 594 1072
rect 622 1068 626 1072
rect 70 1058 74 1062
rect 94 1059 98 1063
rect 158 1058 162 1062
rect 230 1058 234 1062
rect 254 1059 258 1063
rect 286 1058 290 1062
rect 406 1058 410 1062
rect 438 1058 442 1062
rect 470 1058 474 1062
rect 502 1058 506 1062
rect 582 1058 586 1062
rect 622 1058 626 1062
rect 654 1068 658 1072
rect 670 1068 674 1072
rect 878 1068 882 1072
rect 990 1068 994 1072
rect 1166 1068 1170 1072
rect 1214 1068 1218 1072
rect 1254 1078 1258 1082
rect 1278 1068 1282 1072
rect 1318 1068 1322 1072
rect 1342 1078 1346 1082
rect 1382 1078 1386 1082
rect 1398 1068 1402 1072
rect 726 1058 730 1062
rect 782 1058 786 1062
rect 806 1058 810 1062
rect 846 1058 850 1062
rect 894 1059 898 1063
rect 1014 1058 1018 1062
rect 1094 1058 1098 1062
rect 1102 1058 1106 1062
rect 1158 1058 1162 1062
rect 1174 1058 1178 1062
rect 1182 1058 1186 1062
rect 1206 1058 1210 1062
rect 1222 1058 1226 1062
rect 1270 1058 1274 1062
rect 1286 1058 1290 1062
rect 1310 1058 1314 1062
rect 1358 1058 1362 1062
rect 1382 1058 1386 1062
rect 1422 1058 1426 1062
rect 454 1048 458 1052
rect 558 1048 562 1052
rect 598 1048 602 1052
rect 630 1048 634 1052
rect 670 1048 674 1052
rect 1142 1048 1146 1052
rect 1302 1048 1306 1052
rect 654 1038 658 1042
rect 742 1038 746 1042
rect 1286 1038 1290 1042
rect 1110 1018 1114 1022
rect 1190 1018 1194 1022
rect 472 1003 476 1007
rect 477 1003 481 1007
rect 482 1003 486 1007
rect 446 988 450 992
rect 550 988 554 992
rect 614 988 618 992
rect 814 988 818 992
rect 894 988 898 992
rect 950 988 954 992
rect 966 988 970 992
rect 998 988 1002 992
rect 1486 988 1490 992
rect 6 978 10 982
rect 1422 978 1426 982
rect 30 968 34 972
rect 70 968 74 972
rect 150 968 154 972
rect 582 968 586 972
rect 646 968 650 972
rect 1254 968 1258 972
rect 1366 968 1370 972
rect 326 958 330 962
rect 566 958 570 962
rect 654 958 658 962
rect 1118 958 1122 962
rect 1150 958 1154 962
rect 1166 958 1170 962
rect 1238 958 1242 962
rect 1270 958 1274 962
rect 22 948 26 952
rect 118 947 122 951
rect 214 947 218 951
rect 262 948 266 952
rect 310 948 314 952
rect 334 948 338 952
rect 350 948 354 952
rect 406 948 410 952
rect 414 948 418 952
rect 446 948 450 952
rect 510 948 514 952
rect 542 948 546 952
rect 574 948 578 952
rect 598 948 602 952
rect 622 948 626 952
rect 678 948 682 952
rect 702 948 706 952
rect 718 948 722 952
rect 750 947 754 951
rect 782 948 786 952
rect 822 948 826 952
rect 862 948 866 952
rect 878 948 882 952
rect 902 948 906 952
rect 910 948 914 952
rect 918 948 922 952
rect 1054 948 1058 952
rect 1086 947 1090 951
rect 1134 948 1138 952
rect 1174 948 1178 952
rect 1190 948 1194 952
rect 1222 948 1226 952
rect 1254 948 1258 952
rect 62 938 66 942
rect 94 938 98 942
rect 134 938 138 942
rect 230 938 234 942
rect 246 938 250 942
rect 294 938 298 942
rect 302 938 306 942
rect 318 938 322 942
rect 358 938 362 942
rect 406 938 410 942
rect 502 938 506 942
rect 534 938 538 942
rect 574 938 578 942
rect 630 938 634 942
rect 678 938 682 942
rect 974 938 978 942
rect 1126 938 1130 942
rect 1142 938 1146 942
rect 1174 938 1178 942
rect 1302 947 1306 951
rect 1334 948 1338 952
rect 1398 948 1402 952
rect 1406 948 1410 952
rect 1446 948 1450 952
rect 1246 938 1250 942
rect 1374 938 1378 942
rect 1390 938 1394 942
rect 1430 938 1434 942
rect 182 928 186 932
rect 334 928 338 932
rect 430 928 434 932
rect 486 928 490 932
rect 518 928 522 932
rect 526 928 530 932
rect 558 928 562 932
rect 686 928 690 932
rect 942 928 946 932
rect 1038 928 1042 932
rect 1374 928 1378 932
rect 1438 928 1442 932
rect 374 918 378 922
rect 950 918 954 922
rect 1238 918 1242 922
rect 976 903 980 907
rect 981 903 985 907
rect 986 903 990 907
rect 142 888 146 892
rect 230 888 234 892
rect 270 888 274 892
rect 430 888 434 892
rect 518 888 522 892
rect 582 888 586 892
rect 614 888 618 892
rect 702 888 706 892
rect 758 888 762 892
rect 894 888 898 892
rect 966 888 970 892
rect 1030 888 1034 892
rect 1142 888 1146 892
rect 1214 888 1218 892
rect 1430 888 1434 892
rect 46 878 50 882
rect 94 878 98 882
rect 246 878 250 882
rect 278 878 282 882
rect 566 878 570 882
rect 654 878 658 882
rect 6 868 10 872
rect 126 868 130 872
rect 174 868 178 872
rect 182 868 186 872
rect 286 868 290 872
rect 334 868 338 872
rect 350 868 354 872
rect 478 868 482 872
rect 510 868 514 872
rect 542 868 546 872
rect 558 868 562 872
rect 566 868 570 872
rect 638 868 642 872
rect 662 868 666 872
rect 726 868 730 872
rect 774 868 778 872
rect 862 868 866 872
rect 958 868 962 872
rect 990 868 994 872
rect 1038 868 1042 872
rect 1070 868 1074 872
rect 1102 868 1106 872
rect 1166 868 1170 872
rect 1206 868 1210 872
rect 1334 868 1338 872
rect 1486 868 1490 872
rect 94 859 98 863
rect 190 858 194 862
rect 214 858 218 862
rect 374 858 378 862
rect 454 858 458 862
rect 502 858 506 862
rect 510 858 514 862
rect 534 858 538 862
rect 542 858 546 862
rect 574 858 578 862
rect 590 858 594 862
rect 630 858 634 862
rect 654 858 658 862
rect 694 858 698 862
rect 718 858 722 862
rect 838 858 842 862
rect 878 858 882 862
rect 934 858 938 862
rect 982 858 986 862
rect 1014 858 1018 862
rect 1078 858 1082 862
rect 1110 858 1114 862
rect 1142 858 1146 862
rect 1158 858 1162 862
rect 1190 858 1194 862
rect 1294 859 1298 863
rect 1350 859 1354 863
rect 1446 858 1450 862
rect 1454 858 1458 862
rect 206 848 210 852
rect 462 848 466 852
rect 478 848 482 852
rect 518 848 522 852
rect 606 848 610 852
rect 638 848 642 852
rect 686 848 690 852
rect 966 848 970 852
rect 1084 848 1088 852
rect 1094 848 1098 852
rect 1198 848 1202 852
rect 302 838 306 842
rect 446 838 450 842
rect 590 838 594 842
rect 782 838 786 842
rect 798 838 802 842
rect 1182 838 1186 842
rect 1414 838 1418 842
rect 454 828 458 832
rect 190 818 194 822
rect 1190 818 1194 822
rect 1230 818 1234 822
rect 1430 818 1434 822
rect 472 803 476 807
rect 477 803 481 807
rect 482 803 486 807
rect 182 788 186 792
rect 278 788 282 792
rect 342 788 346 792
rect 438 788 442 792
rect 534 788 538 792
rect 614 788 618 792
rect 742 788 746 792
rect 870 788 874 792
rect 934 788 938 792
rect 966 788 970 792
rect 1302 788 1306 792
rect 1486 788 1490 792
rect 894 778 898 782
rect 6 768 10 772
rect 158 768 162 772
rect 862 768 866 772
rect 886 768 890 772
rect 974 768 978 772
rect 1078 768 1082 772
rect 1086 768 1090 772
rect 1142 768 1146 772
rect 1382 768 1386 772
rect 126 758 130 762
rect 174 758 178 762
rect 206 758 210 762
rect 262 758 266 762
rect 390 758 394 762
rect 406 758 410 762
rect 470 758 474 762
rect 494 758 498 762
rect 806 758 810 762
rect 814 758 818 762
rect 846 758 850 762
rect 902 758 906 762
rect 958 758 962 762
rect 990 758 994 762
rect 1094 758 1098 762
rect 1126 758 1130 762
rect 1158 758 1162 762
rect 1244 758 1248 762
rect 1254 758 1258 762
rect 1318 758 1322 762
rect 1366 758 1370 762
rect 38 748 42 752
rect 62 748 66 752
rect 134 748 138 752
rect 190 748 194 752
rect 294 748 298 752
rect 310 748 314 752
rect 382 748 386 752
rect 430 748 434 752
rect 510 748 514 752
rect 70 738 74 742
rect 94 738 98 742
rect 102 740 106 744
rect 678 747 682 751
rect 766 748 770 752
rect 830 748 834 752
rect 854 748 858 752
rect 894 748 898 752
rect 910 748 914 752
rect 918 748 922 752
rect 942 748 946 752
rect 966 748 970 752
rect 1038 748 1042 752
rect 1086 748 1090 752
rect 1118 748 1122 752
rect 1142 748 1146 752
rect 1190 748 1194 752
rect 1206 748 1210 752
rect 1230 748 1234 752
rect 1270 748 1274 752
rect 1302 748 1306 752
rect 1350 748 1354 752
rect 1382 748 1386 752
rect 1430 748 1434 752
rect 1438 748 1442 752
rect 126 738 130 742
rect 158 738 162 742
rect 230 738 234 742
rect 246 738 250 742
rect 366 738 370 742
rect 406 738 410 742
rect 430 738 434 742
rect 454 738 458 742
rect 510 738 514 742
rect 518 738 522 742
rect 558 738 562 742
rect 566 738 570 742
rect 574 738 578 742
rect 694 738 698 742
rect 710 738 714 742
rect 790 738 794 742
rect 838 738 842 742
rect 1046 738 1050 742
rect 1062 738 1066 742
rect 1102 738 1106 742
rect 1134 738 1138 742
rect 1182 738 1186 742
rect 1198 738 1202 742
rect 1230 738 1234 742
rect 1262 738 1266 742
rect 1326 738 1330 742
rect 1342 738 1346 742
rect 1422 738 1426 742
rect 62 728 66 732
rect 238 728 242 732
rect 278 728 282 732
rect 302 728 306 732
rect 326 728 330 732
rect 374 728 378 732
rect 398 728 402 732
rect 446 728 450 732
rect 494 728 498 732
rect 542 728 546 732
rect 782 728 786 732
rect 1054 728 1058 732
rect 1166 728 1170 732
rect 1406 728 1410 732
rect 70 718 74 722
rect 174 718 178 722
rect 262 718 266 722
rect 478 718 482 722
rect 550 718 554 722
rect 798 718 802 722
rect 1174 718 1178 722
rect 1222 718 1226 722
rect 1334 718 1338 722
rect 976 703 980 707
rect 981 703 985 707
rect 986 703 990 707
rect 406 688 410 692
rect 542 688 546 692
rect 678 688 682 692
rect 726 688 730 692
rect 782 688 786 692
rect 814 688 818 692
rect 830 688 834 692
rect 878 688 882 692
rect 998 688 1002 692
rect 1150 688 1154 692
rect 1294 688 1298 692
rect 1390 688 1394 692
rect 1486 688 1490 692
rect 214 678 218 682
rect 398 678 402 682
rect 454 678 458 682
rect 550 678 554 682
rect 790 678 794 682
rect 822 678 826 682
rect 910 678 914 682
rect 942 678 946 682
rect 1006 678 1010 682
rect 1166 678 1170 682
rect 1246 678 1250 682
rect 1302 678 1306 682
rect 1406 678 1410 682
rect 1446 678 1450 682
rect 6 668 10 672
rect 46 668 50 672
rect 110 668 114 672
rect 126 668 130 672
rect 190 668 194 672
rect 206 668 210 672
rect 254 668 258 672
rect 318 668 322 672
rect 382 668 386 672
rect 422 668 426 672
rect 430 668 434 672
rect 470 668 474 672
rect 542 668 546 672
rect 558 668 562 672
rect 614 668 618 672
rect 654 668 658 672
rect 702 668 706 672
rect 806 668 810 672
rect 854 668 858 672
rect 862 668 866 672
rect 886 668 890 672
rect 926 668 930 672
rect 1046 668 1050 672
rect 1062 668 1066 672
rect 1102 668 1106 672
rect 1126 668 1130 672
rect 1222 668 1226 672
rect 1262 668 1266 672
rect 1270 668 1274 672
rect 1318 668 1322 672
rect 1358 668 1362 672
rect 1366 668 1370 672
rect 1398 668 1402 672
rect 1406 668 1410 672
rect 94 659 98 663
rect 142 658 146 662
rect 158 658 162 662
rect 198 658 202 662
rect 246 658 250 662
rect 278 658 282 662
rect 310 658 314 662
rect 334 658 338 662
rect 374 658 378 662
rect 486 658 490 662
rect 534 658 538 662
rect 550 658 554 662
rect 566 658 570 662
rect 646 658 650 662
rect 702 658 706 662
rect 774 658 778 662
rect 806 658 810 662
rect 846 658 850 662
rect 910 658 914 662
rect 926 658 930 662
rect 958 658 962 662
rect 1030 658 1034 662
rect 1046 658 1050 662
rect 1086 658 1090 662
rect 1110 658 1114 662
rect 1150 658 1154 662
rect 1182 658 1186 662
rect 1198 658 1202 662
rect 1230 658 1234 662
rect 1262 658 1266 662
rect 1278 658 1282 662
rect 1326 658 1330 662
rect 1358 658 1362 662
rect 1374 658 1378 662
rect 1414 658 1418 662
rect 1454 658 1458 662
rect 230 648 234 652
rect 286 648 290 652
rect 326 648 330 652
rect 358 648 362 652
rect 374 648 378 652
rect 406 648 410 652
rect 590 648 594 652
rect 614 648 618 652
rect 630 648 634 652
rect 878 648 882 652
rect 902 648 906 652
rect 1038 648 1042 652
rect 1094 648 1098 652
rect 1126 648 1130 652
rect 1158 648 1162 652
rect 1174 648 1178 652
rect 1190 648 1194 652
rect 1246 648 1250 652
rect 1294 648 1298 652
rect 1344 648 1348 652
rect 1390 648 1394 652
rect 1430 648 1434 652
rect 270 638 274 642
rect 342 638 346 642
rect 350 638 354 642
rect 1062 638 1066 642
rect 1078 638 1082 642
rect 1142 638 1146 642
rect 1334 638 1338 642
rect 1198 628 1202 632
rect 310 618 314 622
rect 438 618 442 622
rect 1302 618 1306 622
rect 1438 618 1442 622
rect 472 603 476 607
rect 477 603 481 607
rect 482 603 486 607
rect 94 588 98 592
rect 966 588 970 592
rect 1102 588 1106 592
rect 1190 588 1194 592
rect 1334 588 1338 592
rect 1462 588 1466 592
rect 6 578 10 582
rect 334 578 338 582
rect 878 578 882 582
rect 1446 578 1450 582
rect 30 568 34 572
rect 110 568 114 572
rect 1134 568 1138 572
rect 1254 568 1258 572
rect 1294 568 1298 572
rect 1398 568 1402 572
rect 1422 568 1426 572
rect 1478 568 1482 572
rect 398 558 402 562
rect 582 558 586 562
rect 726 558 730 562
rect 22 548 26 552
rect 46 548 50 552
rect 86 548 90 552
rect 158 547 162 551
rect 222 548 226 552
rect 270 547 274 551
rect 342 548 346 552
rect 390 548 394 552
rect 542 548 546 552
rect 630 548 634 552
rect 702 548 706 552
rect 750 548 754 552
rect 806 548 810 552
rect 814 548 818 552
rect 846 558 850 562
rect 1118 558 1122 562
rect 910 548 914 552
rect 926 548 930 552
rect 942 548 946 552
rect 1030 547 1034 551
rect 1062 548 1066 552
rect 1086 548 1090 552
rect 1134 548 1138 552
rect 1158 548 1162 552
rect 1190 548 1194 552
rect 1214 558 1218 562
rect 1238 548 1242 552
rect 1254 548 1258 552
rect 1302 548 1306 552
rect 1358 548 1362 552
rect 1374 548 1378 552
rect 1422 548 1426 552
rect 174 538 178 542
rect 190 538 194 542
rect 238 538 242 542
rect 254 538 258 542
rect 366 538 370 542
rect 414 538 418 542
rect 422 538 426 542
rect 470 538 474 542
rect 494 538 498 542
rect 542 538 546 542
rect 598 540 602 544
rect 646 538 650 542
rect 670 538 674 542
rect 678 538 682 542
rect 710 538 714 542
rect 750 538 754 542
rect 782 538 786 542
rect 814 538 818 542
rect 870 538 874 542
rect 918 538 922 542
rect 934 538 938 542
rect 1046 538 1050 542
rect 1142 538 1146 542
rect 1238 538 1242 542
rect 1246 538 1250 542
rect 1278 538 1282 542
rect 1310 538 1314 542
rect 1406 538 1410 542
rect 1454 538 1458 542
rect 54 528 58 532
rect 406 528 410 532
rect 614 528 618 532
rect 646 528 650 532
rect 662 528 666 532
rect 758 528 762 532
rect 774 528 778 532
rect 870 528 874 532
rect 902 528 906 532
rect 1078 528 1082 532
rect 1326 528 1330 532
rect 1374 528 1378 532
rect 62 518 66 522
rect 446 518 450 522
rect 510 518 514 522
rect 566 518 570 522
rect 742 518 746 522
rect 838 518 842 522
rect 894 518 898 522
rect 1070 518 1074 522
rect 1318 518 1322 522
rect 1414 518 1418 522
rect 976 503 980 507
rect 981 503 985 507
rect 986 503 990 507
rect 6 488 10 492
rect 366 488 370 492
rect 798 488 802 492
rect 830 488 834 492
rect 1134 488 1138 492
rect 1262 488 1266 492
rect 1454 488 1458 492
rect 102 478 106 482
rect 254 478 258 482
rect 550 478 554 482
rect 622 478 626 482
rect 662 478 666 482
rect 726 478 730 482
rect 734 478 738 482
rect 750 478 754 482
rect 774 478 778 482
rect 822 478 826 482
rect 1022 478 1026 482
rect 86 468 90 472
rect 174 468 178 472
rect 246 468 250 472
rect 254 468 258 472
rect 302 468 306 472
rect 638 468 642 472
rect 670 468 674 472
rect 694 468 698 472
rect 710 468 714 472
rect 814 468 818 472
rect 862 468 866 472
rect 894 468 898 472
rect 910 468 914 472
rect 926 468 930 472
rect 1078 468 1082 472
rect 1126 468 1130 472
rect 1182 468 1186 472
rect 1278 468 1282 472
rect 1286 468 1290 472
rect 1302 478 1306 482
rect 1358 478 1362 482
rect 1470 478 1474 482
rect 1350 468 1354 472
rect 1390 468 1394 472
rect 1422 468 1426 472
rect 70 459 74 463
rect 102 458 106 462
rect 118 458 122 462
rect 126 458 130 462
rect 166 458 170 462
rect 198 458 202 462
rect 206 458 210 462
rect 286 458 290 462
rect 310 458 314 462
rect 342 458 346 462
rect 430 459 434 463
rect 510 458 514 462
rect 534 458 538 462
rect 574 458 578 462
rect 598 458 602 462
rect 750 458 754 462
rect 758 458 762 462
rect 838 458 842 462
rect 886 458 890 462
rect 902 458 906 462
rect 934 458 938 462
rect 958 458 962 462
rect 966 458 970 462
rect 1006 458 1010 462
rect 1086 458 1090 462
rect 1142 458 1146 462
rect 1214 458 1218 462
rect 1270 458 1274 462
rect 1318 458 1322 462
rect 1342 458 1346 462
rect 1382 458 1386 462
rect 1406 458 1410 462
rect 1446 458 1450 462
rect 302 448 306 452
rect 342 448 346 452
rect 686 448 690 452
rect 806 448 810 452
rect 846 448 850 452
rect 942 448 946 452
rect 1326 448 1330 452
rect 1398 448 1402 452
rect 254 438 258 442
rect 278 438 282 442
rect 566 438 570 442
rect 886 438 890 442
rect 926 438 930 442
rect 958 438 962 442
rect 1046 438 1050 442
rect 238 418 242 422
rect 286 418 290 422
rect 358 418 362 422
rect 590 418 594 422
rect 614 418 618 422
rect 1030 418 1034 422
rect 1158 418 1162 422
rect 1342 418 1346 422
rect 1366 418 1370 422
rect 472 403 476 407
rect 477 403 481 407
rect 482 403 486 407
rect 230 388 234 392
rect 758 388 762 392
rect 1206 388 1210 392
rect 1334 388 1338 392
rect 1398 388 1402 392
rect 1430 378 1434 382
rect 6 368 10 372
rect 222 368 226 372
rect 254 368 258 372
rect 766 368 770 372
rect 1486 368 1490 372
rect 182 358 186 362
rect 190 358 194 362
rect 238 358 242 362
rect 388 358 392 362
rect 398 358 402 362
rect 406 358 410 362
rect 454 358 458 362
rect 462 358 466 362
rect 526 358 530 362
rect 582 358 586 362
rect 654 358 658 362
rect 726 358 730 362
rect 750 358 754 362
rect 854 358 858 362
rect 1036 358 1040 362
rect 1054 358 1058 362
rect 1110 358 1114 362
rect 94 347 98 351
rect 158 348 162 352
rect 230 348 234 352
rect 278 348 282 352
rect 294 348 298 352
rect 310 348 314 352
rect 326 348 330 352
rect 334 348 338 352
rect 374 348 378 352
rect 510 348 514 352
rect 518 348 522 352
rect 526 348 530 352
rect 574 348 578 352
rect 598 348 602 352
rect 614 348 618 352
rect 686 348 690 352
rect 758 348 762 352
rect 798 348 802 352
rect 846 348 850 352
rect 878 348 882 352
rect 902 348 906 352
rect 982 348 986 352
rect 1014 348 1018 352
rect 1030 348 1034 352
rect 1062 348 1066 352
rect 1094 348 1098 352
rect 1102 348 1106 352
rect 86 338 90 342
rect 142 338 146 342
rect 166 338 170 342
rect 206 338 210 342
rect 286 338 290 342
rect 374 338 378 342
rect 422 338 426 342
rect 438 338 442 342
rect 518 338 522 342
rect 550 338 554 342
rect 606 338 610 342
rect 630 338 634 342
rect 638 338 642 342
rect 742 338 746 342
rect 918 338 922 342
rect 942 338 946 342
rect 990 338 994 342
rect 1022 338 1026 342
rect 1054 338 1058 342
rect 1142 347 1146 351
rect 1214 348 1218 352
rect 1278 348 1282 352
rect 1342 348 1346 352
rect 1374 348 1378 352
rect 1414 348 1418 352
rect 1438 348 1442 352
rect 1126 338 1130 342
rect 1222 338 1226 342
rect 1254 338 1258 342
rect 1350 338 1354 342
rect 62 328 66 332
rect 126 328 130 332
rect 310 328 314 332
rect 334 328 338 332
rect 366 328 370 332
rect 430 328 434 332
rect 462 328 466 332
rect 558 328 562 332
rect 670 328 674 332
rect 830 328 834 332
rect 894 328 898 332
rect 934 328 938 332
rect 1238 328 1242 332
rect 1390 328 1394 332
rect 1406 328 1410 332
rect 174 318 178 322
rect 190 318 194 322
rect 358 318 362 322
rect 446 318 450 322
rect 582 318 586 322
rect 662 318 666 322
rect 694 318 698 322
rect 710 318 714 322
rect 814 318 818 322
rect 1230 318 1234 322
rect 1334 318 1338 322
rect 1358 318 1362 322
rect 976 303 980 307
rect 981 303 985 307
rect 986 303 990 307
rect 6 288 10 292
rect 198 288 202 292
rect 262 288 266 292
rect 878 288 882 292
rect 982 288 986 292
rect 1270 288 1274 292
rect 1286 288 1290 292
rect 1318 288 1322 292
rect 1446 288 1450 292
rect 206 278 210 282
rect 270 278 274 282
rect 358 278 362 282
rect 390 278 394 282
rect 454 278 458 282
rect 534 278 538 282
rect 622 278 626 282
rect 662 278 666 282
rect 790 278 794 282
rect 1142 278 1146 282
rect 1294 278 1298 282
rect 1350 278 1354 282
rect 86 268 90 272
rect 166 268 170 272
rect 206 268 210 272
rect 222 268 226 272
rect 238 268 242 272
rect 318 268 322 272
rect 366 268 370 272
rect 390 268 394 272
rect 398 268 402 272
rect 414 268 418 272
rect 438 268 442 272
rect 478 268 482 272
rect 518 268 522 272
rect 534 268 538 272
rect 598 268 602 272
rect 678 268 682 272
rect 718 268 722 272
rect 766 268 770 272
rect 798 268 802 272
rect 862 268 866 272
rect 870 268 874 272
rect 1158 268 1162 272
rect 1190 268 1194 272
rect 1310 268 1314 272
rect 1366 268 1370 272
rect 1382 268 1386 272
rect 1486 268 1490 272
rect 70 259 74 263
rect 118 258 122 262
rect 198 258 202 262
rect 230 258 234 262
rect 254 258 258 262
rect 310 258 314 262
rect 318 258 322 262
rect 366 258 370 262
rect 406 258 410 262
rect 422 258 426 262
rect 454 258 458 262
rect 486 258 490 262
rect 510 258 514 262
rect 518 258 522 262
rect 534 258 538 262
rect 558 258 562 262
rect 574 258 578 262
rect 590 258 594 262
rect 606 258 610 262
rect 646 258 650 262
rect 686 258 690 262
rect 726 258 730 262
rect 758 258 762 262
rect 766 258 770 262
rect 806 258 810 262
rect 918 258 922 262
rect 942 258 946 262
rect 982 258 986 262
rect 1022 258 1026 262
rect 1078 258 1082 262
rect 1110 259 1114 263
rect 1174 258 1178 262
rect 1230 258 1234 262
rect 1278 258 1282 262
rect 1302 258 1306 262
rect 1334 258 1338 262
rect 1390 258 1394 262
rect 1454 258 1458 262
rect 102 248 106 252
rect 134 248 138 252
rect 246 248 250 252
rect 502 248 506 252
rect 566 248 570 252
rect 614 248 618 252
rect 654 248 658 252
rect 758 248 762 252
rect 822 248 826 252
rect 846 248 850 252
rect 550 238 554 242
rect 566 238 570 242
rect 638 238 642 242
rect 1046 238 1050 242
rect 118 218 122 222
rect 286 218 290 222
rect 646 218 650 222
rect 710 218 714 222
rect 774 218 778 222
rect 830 218 834 222
rect 878 218 882 222
rect 1014 218 1018 222
rect 1038 218 1042 222
rect 472 203 476 207
rect 477 203 481 207
rect 482 203 486 207
rect 62 188 66 192
rect 102 188 106 192
rect 230 188 234 192
rect 254 188 258 192
rect 310 188 314 192
rect 550 188 554 192
rect 614 188 618 192
rect 646 188 650 192
rect 1462 188 1466 192
rect 694 178 698 182
rect 206 168 210 172
rect 262 168 266 172
rect 422 168 426 172
rect 430 168 434 172
rect 1246 168 1250 172
rect 222 158 226 162
rect 238 158 242 162
rect 286 158 290 162
rect 318 158 322 162
rect 326 158 330 162
rect 390 158 394 162
rect 414 158 418 162
rect 534 158 538 162
rect 574 158 578 162
rect 654 158 658 162
rect 966 158 970 162
rect 62 148 66 152
rect 134 148 138 152
rect 166 147 170 151
rect 198 148 202 152
rect 214 148 218 152
rect 254 148 258 152
rect 294 148 298 152
rect 318 148 322 152
rect 358 148 362 152
rect 430 148 434 152
rect 454 148 458 152
rect 518 148 522 152
rect 558 148 562 152
rect 662 148 666 152
rect 686 148 690 152
rect 726 148 730 152
rect 774 148 778 152
rect 814 148 818 152
rect 878 148 882 152
rect 910 148 914 152
rect 942 148 946 152
rect 1006 148 1010 152
rect 1054 148 1058 152
rect 1078 148 1082 152
rect 1110 148 1114 152
rect 1150 148 1154 152
rect 1206 148 1210 152
rect 1214 148 1218 152
rect 1294 148 1298 152
rect 86 138 90 142
rect 302 138 306 142
rect 350 138 354 142
rect 374 138 378 142
rect 414 138 418 142
rect 454 138 458 142
rect 494 138 498 142
rect 526 138 530 142
rect 558 138 562 142
rect 566 138 570 142
rect 590 138 594 142
rect 638 138 642 142
rect 1374 147 1378 151
rect 1446 148 1450 152
rect 718 138 722 142
rect 742 138 746 142
rect 806 138 810 142
rect 846 138 850 142
rect 958 138 962 142
rect 982 138 986 142
rect 1014 138 1018 142
rect 1086 138 1090 142
rect 1102 138 1106 142
rect 1174 138 1178 142
rect 1230 138 1234 142
rect 1382 138 1386 142
rect 238 128 242 132
rect 278 128 282 132
rect 358 128 362 132
rect 390 128 394 132
rect 470 128 474 132
rect 518 128 522 132
rect 606 128 610 132
rect 630 128 634 132
rect 678 128 682 132
rect 710 128 714 132
rect 750 128 754 132
rect 790 128 794 132
rect 854 128 858 132
rect 934 128 938 132
rect 1038 128 1042 132
rect 1062 128 1066 132
rect 1246 128 1250 132
rect 6 118 10 122
rect 366 118 370 122
rect 438 118 442 122
rect 742 118 746 122
rect 806 118 810 122
rect 870 118 874 122
rect 926 118 930 122
rect 950 118 954 122
rect 1022 118 1026 122
rect 1190 118 1194 122
rect 1438 118 1442 122
rect 1462 118 1466 122
rect 976 103 980 107
rect 981 103 985 107
rect 986 103 990 107
rect 62 88 66 92
rect 166 88 170 92
rect 270 88 274 92
rect 374 88 378 92
rect 430 88 434 92
rect 558 88 562 92
rect 702 88 706 92
rect 934 88 938 92
rect 1302 88 1306 92
rect 1454 88 1458 92
rect 70 78 74 82
rect 78 78 82 82
rect 166 78 170 82
rect 206 78 210 82
rect 222 78 226 82
rect 366 78 370 82
rect 470 78 474 82
rect 534 78 538 82
rect 1070 78 1074 82
rect 6 68 10 72
rect 30 68 34 72
rect 46 68 50 72
rect 54 68 58 72
rect 78 68 82 72
rect 102 68 106 72
rect 118 68 122 72
rect 182 68 186 72
rect 230 68 234 72
rect 278 68 282 72
rect 294 68 298 72
rect 350 68 354 72
rect 494 68 498 72
rect 534 68 538 72
rect 590 68 594 72
rect 622 68 626 72
rect 638 68 642 72
rect 782 68 786 72
rect 1270 68 1274 72
rect 1318 68 1322 72
rect 1446 68 1450 72
rect 22 58 26 62
rect 94 58 98 62
rect 158 58 162 62
rect 190 58 194 62
rect 238 58 242 62
rect 302 58 306 62
rect 382 58 386 62
rect 430 58 434 62
rect 462 58 466 62
rect 470 58 474 62
rect 526 58 530 62
rect 550 58 554 62
rect 582 58 586 62
rect 638 58 642 62
rect 646 58 650 62
rect 678 58 682 62
rect 694 58 698 62
rect 758 58 762 62
rect 814 58 818 62
rect 838 58 842 62
rect 878 58 882 62
rect 902 58 906 62
rect 966 58 970 62
rect 1046 58 1050 62
rect 1070 59 1074 63
rect 1102 58 1106 62
rect 1126 58 1130 62
rect 1150 58 1154 62
rect 1174 58 1178 62
rect 1198 58 1202 62
rect 1222 58 1226 62
rect 1246 58 1250 62
rect 1374 58 1378 62
rect 1398 58 1402 62
rect 1422 58 1426 62
rect 102 48 106 52
rect 308 48 312 52
rect 326 48 330 52
rect 422 48 426 52
rect 508 48 512 52
rect 614 48 618 52
rect 622 48 626 52
rect 670 48 674 52
rect 1486 48 1490 52
rect 190 38 194 42
rect 438 38 442 42
rect 686 38 690 42
rect 1006 38 1010 42
rect 662 18 666 22
rect 798 18 802 22
rect 822 18 826 22
rect 958 18 962 22
rect 982 18 986 22
rect 1118 18 1122 22
rect 1142 18 1146 22
rect 1214 18 1218 22
rect 1262 18 1266 22
rect 1342 18 1346 22
rect 1390 18 1394 22
rect 1414 18 1418 22
rect 1438 18 1442 22
rect 472 3 476 7
rect 477 3 481 7
rect 482 3 486 7
<< metal2 >>
rect 102 1192 105 1231
rect 166 1212 169 1231
rect 214 1192 217 1231
rect 478 1228 497 1231
rect 476 1203 477 1207
rect 481 1203 482 1207
rect 486 1203 488 1207
rect 494 1192 497 1228
rect 614 1212 617 1231
rect 702 1192 705 1231
rect 822 1192 825 1231
rect 846 1192 849 1231
rect 862 1228 873 1231
rect 886 1228 897 1231
rect 218 1168 222 1171
rect 6 1132 9 1168
rect 70 1151 73 1158
rect 142 1152 145 1158
rect 198 1152 201 1168
rect 174 1142 177 1148
rect 126 1132 129 1138
rect 178 1128 182 1131
rect 62 1072 65 1078
rect 6 1062 9 1068
rect 70 1062 73 1128
rect 190 1122 193 1128
rect 166 1092 169 1108
rect 254 1082 257 1148
rect 286 1112 289 1147
rect 318 1142 321 1168
rect 662 1162 665 1168
rect 402 1158 406 1161
rect 650 1158 654 1161
rect 394 1148 398 1151
rect 382 1142 385 1148
rect 366 1132 369 1138
rect 334 1112 337 1118
rect 374 1112 377 1138
rect 382 1092 385 1138
rect 406 1122 409 1148
rect 414 1142 417 1148
rect 422 1092 425 1158
rect 638 1152 641 1158
rect 530 1148 534 1151
rect 438 1142 441 1148
rect 454 1132 457 1138
rect 442 1128 446 1131
rect 430 1112 433 1128
rect 394 1078 398 1081
rect 126 1072 129 1078
rect 286 1072 289 1078
rect 202 1068 206 1071
rect 378 1068 382 1071
rect 90 1059 94 1061
rect 142 1062 145 1068
rect 90 1058 97 1059
rect 6 982 9 988
rect 70 972 73 1058
rect 146 968 150 971
rect 22 952 25 968
rect 30 962 33 968
rect 46 882 49 888
rect 62 872 65 938
rect 94 882 97 938
rect 118 922 121 947
rect 134 942 137 948
rect 142 892 145 918
rect 158 902 161 1058
rect 182 932 185 938
rect 126 872 129 878
rect 6 862 9 868
rect 6 762 9 768
rect 62 752 65 868
rect 94 842 97 859
rect 174 851 177 868
rect 182 862 185 868
rect 190 862 193 968
rect 214 951 217 958
rect 230 942 233 1058
rect 254 1052 257 1059
rect 286 1052 289 1058
rect 334 1042 337 1068
rect 398 972 401 1078
rect 414 1062 417 1068
rect 430 1062 433 1108
rect 462 1082 465 1148
rect 646 1142 649 1158
rect 734 1151 737 1158
rect 510 1072 513 1078
rect 518 1072 521 1118
rect 526 1082 529 1118
rect 542 1112 545 1138
rect 550 1122 553 1128
rect 558 1092 561 1128
rect 582 1122 585 1128
rect 598 1092 601 1118
rect 630 1092 633 1108
rect 554 1068 558 1071
rect 586 1068 590 1071
rect 618 1068 622 1071
rect 470 1062 473 1068
rect 502 1062 505 1068
rect 586 1058 590 1061
rect 246 942 249 968
rect 322 958 326 961
rect 262 952 265 958
rect 406 952 409 1058
rect 438 1052 441 1058
rect 454 1052 457 1058
rect 314 948 318 951
rect 330 948 334 951
rect 354 948 358 951
rect 294 942 297 948
rect 322 938 326 941
rect 230 892 233 938
rect 302 922 305 938
rect 358 932 361 938
rect 406 932 409 938
rect 230 872 233 888
rect 246 882 249 908
rect 270 892 273 918
rect 334 912 337 928
rect 414 922 417 948
rect 430 942 433 968
rect 438 962 441 1048
rect 446 992 449 1038
rect 454 952 457 1048
rect 476 1003 477 1007
rect 481 1003 482 1007
rect 486 1003 488 1007
rect 450 948 454 951
rect 502 942 505 1058
rect 550 1048 558 1051
rect 594 1048 598 1051
rect 550 992 553 1048
rect 566 962 569 1048
rect 614 992 617 1038
rect 586 968 590 971
rect 546 948 550 951
rect 494 938 502 941
rect 430 932 433 938
rect 246 862 249 878
rect 218 858 225 861
rect 174 848 185 851
rect 126 762 129 768
rect 134 752 137 828
rect 182 792 185 848
rect 190 832 193 858
rect 210 848 214 851
rect 222 822 225 858
rect 278 852 281 878
rect 286 872 289 888
rect 350 872 353 878
rect 334 862 337 868
rect 374 862 377 918
rect 430 892 433 928
rect 430 862 433 888
rect 450 858 454 861
rect 462 852 465 888
rect 474 868 478 871
rect 486 862 489 928
rect 494 852 497 938
rect 510 931 513 948
rect 526 932 529 938
rect 502 928 513 931
rect 502 862 505 928
rect 518 892 521 928
rect 534 922 537 938
rect 510 872 513 878
rect 534 862 537 888
rect 542 872 545 948
rect 558 932 561 938
rect 566 921 569 958
rect 574 952 577 958
rect 622 952 625 1058
rect 646 1052 649 1118
rect 654 1062 657 1068
rect 634 1048 638 1051
rect 630 962 633 1048
rect 646 962 649 968
rect 654 962 657 1038
rect 574 932 577 938
rect 558 918 569 921
rect 558 872 561 918
rect 582 892 585 918
rect 566 882 569 888
rect 598 882 601 948
rect 622 932 625 948
rect 630 942 633 948
rect 618 888 622 891
rect 650 878 654 881
rect 158 762 161 768
rect 170 758 174 761
rect 190 752 193 818
rect 278 792 281 848
rect 306 838 310 841
rect 442 838 446 841
rect 342 792 345 838
rect 454 832 457 848
rect 478 832 481 848
rect 438 792 441 828
rect 476 803 477 807
rect 481 803 482 807
rect 486 803 488 807
rect 510 782 513 858
rect 518 832 521 848
rect 534 792 537 838
rect 38 732 41 748
rect 70 742 73 748
rect 62 732 65 738
rect 94 732 97 738
rect 58 728 62 731
rect 42 668 46 671
rect 6 662 9 668
rect 62 592 65 728
rect 102 722 105 740
rect 122 738 126 741
rect 158 732 161 738
rect 206 732 209 758
rect 246 742 249 768
rect 258 758 262 761
rect 234 738 238 741
rect 254 732 257 758
rect 310 752 313 758
rect 298 748 302 751
rect 278 732 281 738
rect 242 728 246 731
rect 298 728 302 731
rect 70 692 73 718
rect 126 682 129 718
rect 174 702 177 718
rect 126 672 129 678
rect 190 672 193 678
rect 206 672 209 698
rect 218 678 222 681
rect 94 652 97 659
rect 90 588 94 591
rect 6 582 9 588
rect 110 572 113 668
rect 142 662 145 668
rect 202 658 206 661
rect 158 652 161 658
rect 230 652 233 728
rect 258 718 262 721
rect 254 672 257 688
rect 250 658 254 661
rect 234 648 241 651
rect 30 562 33 568
rect 50 548 54 551
rect 90 548 94 551
rect 158 551 161 558
rect 22 532 25 548
rect 50 528 54 531
rect 6 492 9 528
rect 62 492 65 518
rect 102 482 105 488
rect 86 472 89 478
rect 70 463 73 468
rect 70 458 73 459
rect 6 362 9 368
rect 86 342 89 468
rect 102 462 105 468
rect 118 462 121 468
rect 126 462 129 548
rect 190 542 193 588
rect 238 562 241 648
rect 270 642 273 688
rect 278 662 281 668
rect 286 652 289 728
rect 310 662 313 728
rect 326 722 329 728
rect 318 672 321 718
rect 326 652 329 668
rect 334 662 337 668
rect 358 662 361 778
rect 390 762 393 768
rect 406 762 409 768
rect 466 758 470 761
rect 426 748 430 751
rect 370 738 374 741
rect 370 728 374 731
rect 382 722 385 748
rect 402 738 406 741
rect 458 738 462 741
rect 402 728 409 731
rect 382 672 385 718
rect 406 692 409 728
rect 430 682 433 738
rect 494 732 497 758
rect 510 752 513 778
rect 514 748 518 751
rect 506 738 510 741
rect 450 728 454 731
rect 454 682 457 728
rect 518 722 521 738
rect 542 732 545 858
rect 566 852 569 868
rect 574 862 577 868
rect 586 858 590 861
rect 566 742 569 748
rect 574 742 577 778
rect 554 738 558 741
rect 482 718 486 721
rect 542 692 545 698
rect 550 692 553 718
rect 398 672 401 678
rect 542 672 545 678
rect 418 668 422 671
rect 374 662 377 668
rect 358 652 361 658
rect 406 652 409 658
rect 430 652 433 668
rect 378 648 382 651
rect 350 642 353 648
rect 338 638 342 641
rect 310 592 313 618
rect 338 578 342 581
rect 218 548 222 551
rect 238 542 241 558
rect 390 552 393 618
rect 398 562 401 588
rect 346 548 350 551
rect 174 482 177 538
rect 254 532 257 538
rect 270 522 273 547
rect 174 472 177 478
rect 126 452 129 458
rect 94 351 97 358
rect 62 332 65 338
rect 6 292 9 298
rect 86 272 89 338
rect 126 332 129 338
rect 70 263 73 268
rect 70 258 73 259
rect 62 152 65 188
rect 86 152 89 268
rect 102 252 105 258
rect 118 252 121 258
rect 134 252 137 378
rect 158 352 161 468
rect 166 452 169 458
rect 182 362 185 498
rect 198 462 201 468
rect 206 462 209 468
rect 206 452 209 458
rect 190 362 193 438
rect 230 392 233 518
rect 254 482 257 498
rect 246 472 249 478
rect 238 382 241 418
rect 226 368 230 371
rect 226 348 230 351
rect 142 342 145 348
rect 170 338 174 341
rect 166 272 169 338
rect 106 188 110 191
rect 86 142 89 148
rect 10 118 14 121
rect 6 62 9 68
rect 22 62 25 118
rect 62 92 65 128
rect 70 82 73 88
rect 82 78 86 81
rect 30 72 33 78
rect 42 68 46 71
rect 54 62 57 68
rect 78 62 81 68
rect 94 62 97 108
rect 102 72 105 78
rect 110 61 113 168
rect 118 92 121 218
rect 134 172 137 248
rect 166 192 169 268
rect 174 262 177 318
rect 190 252 193 318
rect 198 292 201 348
rect 210 338 214 341
rect 206 282 209 288
rect 198 262 201 278
rect 238 272 241 358
rect 246 302 249 468
rect 254 462 257 468
rect 286 462 289 478
rect 302 472 305 518
rect 302 452 305 468
rect 310 462 313 498
rect 342 472 345 548
rect 366 542 369 548
rect 366 492 369 508
rect 390 501 393 548
rect 406 542 409 648
rect 470 642 473 668
rect 550 662 553 678
rect 486 652 489 658
rect 534 642 537 658
rect 558 642 561 668
rect 414 542 417 558
rect 438 552 441 618
rect 566 611 569 658
rect 574 652 577 738
rect 566 608 577 611
rect 476 603 477 607
rect 481 603 482 607
rect 486 603 488 607
rect 542 552 545 578
rect 546 548 550 551
rect 422 542 425 548
rect 470 542 473 548
rect 546 538 553 541
rect 402 528 406 531
rect 422 512 425 538
rect 494 532 497 538
rect 390 498 401 501
rect 338 458 342 461
rect 278 442 281 448
rect 258 438 262 441
rect 254 362 257 368
rect 278 352 281 358
rect 286 352 289 418
rect 286 332 289 338
rect 266 288 270 291
rect 206 262 209 268
rect 190 171 193 248
rect 222 211 225 268
rect 230 221 233 258
rect 246 242 249 248
rect 230 218 241 221
rect 222 208 233 211
rect 230 192 233 208
rect 182 168 193 171
rect 206 172 209 178
rect 134 152 137 158
rect 166 151 169 158
rect 166 92 169 118
rect 182 112 185 168
rect 238 162 241 218
rect 254 192 257 258
rect 270 222 273 278
rect 198 152 201 158
rect 222 152 225 158
rect 182 102 185 108
rect 158 82 161 88
rect 162 78 166 81
rect 182 72 185 98
rect 206 82 209 138
rect 214 132 217 148
rect 238 142 241 158
rect 254 152 257 168
rect 262 162 265 168
rect 238 112 241 128
rect 222 82 225 88
rect 122 68 126 71
rect 230 62 233 68
rect 238 62 241 98
rect 102 58 113 61
rect 186 58 190 61
rect 102 52 105 58
rect 158 52 161 58
rect 254 52 257 148
rect 278 132 281 188
rect 286 182 289 218
rect 286 152 289 158
rect 294 152 297 348
rect 302 342 305 448
rect 310 352 313 458
rect 342 442 345 448
rect 358 392 361 418
rect 326 352 329 358
rect 342 352 345 378
rect 398 371 401 498
rect 446 462 449 518
rect 510 462 513 518
rect 550 482 553 538
rect 430 452 433 459
rect 534 422 537 458
rect 566 452 569 518
rect 574 462 577 608
rect 582 572 585 848
rect 590 842 593 848
rect 590 702 593 838
rect 598 772 601 878
rect 662 872 665 1138
rect 678 1132 681 1138
rect 686 1092 689 1148
rect 786 1138 790 1141
rect 750 1112 753 1138
rect 670 1072 673 1078
rect 670 1052 673 1058
rect 678 952 681 1088
rect 742 1082 745 1088
rect 726 1052 729 1058
rect 742 1042 745 1078
rect 782 1062 785 1108
rect 802 1058 806 1061
rect 642 868 646 871
rect 654 862 657 868
rect 634 858 641 861
rect 606 852 609 858
rect 638 852 641 858
rect 654 852 657 858
rect 618 788 622 791
rect 662 752 665 868
rect 678 782 681 938
rect 686 932 689 998
rect 706 948 710 951
rect 750 951 753 958
rect 782 952 785 1058
rect 814 992 817 998
rect 702 892 705 928
rect 718 902 721 948
rect 754 888 758 891
rect 782 882 785 948
rect 822 942 825 948
rect 774 872 777 878
rect 722 868 726 871
rect 778 868 785 871
rect 694 862 697 868
rect 686 842 689 848
rect 718 812 721 858
rect 742 792 745 858
rect 782 842 785 868
rect 822 852 825 938
rect 678 692 681 747
rect 694 742 697 758
rect 710 722 713 738
rect 726 712 729 718
rect 726 692 729 708
rect 766 702 769 748
rect 594 648 598 651
rect 606 651 609 688
rect 702 672 705 678
rect 618 668 622 671
rect 650 668 654 671
rect 774 662 777 778
rect 790 742 793 778
rect 798 762 801 838
rect 830 792 833 1148
rect 846 1002 849 1058
rect 854 942 857 1148
rect 862 1092 865 1228
rect 886 1212 889 1228
rect 910 1212 913 1231
rect 934 1212 937 1231
rect 942 1228 953 1231
rect 870 1192 873 1208
rect 894 1192 897 1208
rect 918 1192 921 1208
rect 942 1192 945 1228
rect 998 1212 1001 1231
rect 1054 1212 1057 1231
rect 1078 1212 1081 1231
rect 1038 1192 1041 1208
rect 1062 1192 1065 1208
rect 1094 1172 1097 1231
rect 1118 1202 1121 1231
rect 874 1148 878 1151
rect 898 1148 902 1151
rect 878 1072 881 1108
rect 926 1092 929 1148
rect 942 1138 950 1141
rect 942 1081 945 1138
rect 978 1118 982 1121
rect 980 1103 981 1107
rect 985 1103 986 1107
rect 990 1103 992 1107
rect 954 1088 958 1091
rect 942 1078 953 1081
rect 926 1072 929 1078
rect 894 992 897 1059
rect 950 992 953 1078
rect 990 1062 993 1068
rect 1014 1062 1017 1118
rect 1022 1102 1025 1148
rect 1046 1112 1049 1148
rect 1074 1138 1078 1141
rect 1086 1112 1089 1118
rect 966 992 969 1048
rect 998 992 1001 1008
rect 902 952 905 968
rect 910 952 913 958
rect 1054 952 1057 1068
rect 862 942 865 948
rect 878 892 881 948
rect 918 942 921 948
rect 894 892 897 938
rect 942 932 945 948
rect 974 932 977 938
rect 838 862 841 888
rect 950 882 953 918
rect 966 892 969 918
rect 980 903 981 907
rect 985 903 986 907
rect 990 903 992 907
rect 1030 892 1033 908
rect 862 872 865 878
rect 1038 872 1041 928
rect 1054 912 1057 948
rect 954 868 958 871
rect 938 858 942 861
rect 870 792 873 828
rect 878 812 881 858
rect 934 792 937 838
rect 942 822 945 858
rect 982 852 985 858
rect 814 762 817 768
rect 786 728 790 731
rect 606 648 614 651
rect 630 642 633 648
rect 582 562 585 568
rect 646 552 649 658
rect 702 552 705 658
rect 774 652 777 658
rect 782 622 785 688
rect 790 672 793 678
rect 698 548 702 551
rect 602 540 606 541
rect 598 538 606 540
rect 614 482 617 528
rect 630 522 633 548
rect 710 542 713 548
rect 642 538 646 541
rect 682 538 686 541
rect 706 538 710 541
rect 658 528 662 531
rect 646 502 649 528
rect 670 482 673 538
rect 626 478 630 481
rect 666 478 670 481
rect 642 468 646 471
rect 598 442 601 458
rect 570 438 574 441
rect 476 403 477 407
rect 481 403 482 407
rect 486 403 488 407
rect 390 368 401 371
rect 390 362 393 368
rect 406 362 409 368
rect 526 362 529 388
rect 392 358 393 362
rect 374 352 377 358
rect 398 352 401 358
rect 338 348 342 351
rect 366 332 369 338
rect 330 328 334 331
rect 310 312 313 328
rect 318 272 321 298
rect 358 291 361 318
rect 374 312 377 338
rect 422 322 425 338
rect 438 332 441 338
rect 454 332 457 358
rect 462 352 465 358
rect 518 352 521 358
rect 530 348 534 351
rect 430 322 433 328
rect 438 311 441 328
rect 430 308 441 311
rect 358 288 369 291
rect 358 272 361 278
rect 366 272 369 288
rect 310 262 313 268
rect 318 251 321 258
rect 310 248 321 251
rect 310 232 313 248
rect 310 192 313 228
rect 326 192 329 238
rect 302 142 305 168
rect 326 162 329 188
rect 314 158 318 161
rect 318 142 321 148
rect 350 142 353 148
rect 358 132 361 148
rect 366 142 369 258
rect 374 251 377 308
rect 390 282 393 288
rect 414 272 417 278
rect 386 268 390 271
rect 398 252 401 268
rect 422 262 425 268
rect 374 248 385 251
rect 374 142 377 148
rect 362 128 366 131
rect 270 92 273 118
rect 366 112 369 118
rect 294 72 297 88
rect 350 72 353 98
rect 382 92 385 248
rect 394 158 398 161
rect 378 88 382 91
rect 362 78 366 81
rect 282 68 286 71
rect 298 58 302 61
rect 326 52 329 58
rect 312 48 313 51
rect 190 42 193 48
rect 310 42 313 48
rect 366 -22 369 78
rect 390 61 393 128
rect 406 112 409 258
rect 430 172 433 308
rect 438 272 441 278
rect 446 272 449 318
rect 454 282 457 328
rect 462 312 465 328
rect 462 302 465 308
rect 510 282 513 348
rect 550 342 553 388
rect 582 362 585 378
rect 578 348 582 351
rect 518 332 521 338
rect 558 332 561 338
rect 574 332 577 348
rect 518 272 521 298
rect 538 278 542 281
rect 538 268 542 271
rect 450 258 454 261
rect 478 242 481 268
rect 574 262 577 268
rect 530 258 534 261
rect 562 258 566 261
rect 582 261 585 318
rect 590 272 593 418
rect 614 372 617 418
rect 610 348 614 351
rect 598 332 601 348
rect 598 322 601 328
rect 606 322 609 338
rect 598 272 601 278
rect 614 271 617 348
rect 630 342 633 378
rect 638 342 641 448
rect 654 362 657 478
rect 678 471 681 538
rect 726 522 729 558
rect 742 548 750 551
rect 742 532 745 548
rect 782 542 785 608
rect 754 538 758 541
rect 762 528 766 531
rect 774 522 777 528
rect 674 468 681 471
rect 694 472 697 498
rect 710 472 713 478
rect 686 452 689 458
rect 654 282 657 358
rect 670 332 673 378
rect 694 352 697 468
rect 686 332 689 348
rect 662 322 665 328
rect 678 322 681 328
rect 710 322 713 328
rect 662 282 665 318
rect 606 268 617 271
rect 582 258 590 261
rect 478 232 481 238
rect 486 232 489 258
rect 502 252 505 258
rect 486 222 489 228
rect 476 203 477 207
rect 481 203 482 207
rect 486 203 488 207
rect 414 142 417 158
rect 422 82 425 168
rect 430 152 433 158
rect 454 152 457 158
rect 454 132 457 138
rect 470 132 473 138
rect 430 92 433 108
rect 438 102 441 118
rect 478 102 481 158
rect 494 142 497 238
rect 510 112 513 258
rect 518 252 521 258
rect 598 252 601 268
rect 606 262 609 268
rect 570 248 577 251
rect 574 242 577 248
rect 554 238 558 241
rect 550 192 553 228
rect 518 152 521 188
rect 526 142 529 178
rect 538 158 542 161
rect 550 141 553 178
rect 558 152 561 168
rect 566 142 569 238
rect 574 162 577 168
rect 550 138 558 141
rect 526 132 529 138
rect 518 122 521 128
rect 470 82 473 88
rect 386 58 393 61
rect 426 58 430 61
rect 438 52 441 68
rect 470 62 473 78
rect 494 72 497 108
rect 490 68 494 71
rect 526 62 529 128
rect 558 92 561 118
rect 566 102 569 138
rect 534 82 537 88
rect 534 62 537 68
rect 550 62 553 78
rect 582 72 585 248
rect 590 172 593 188
rect 606 172 609 258
rect 614 252 617 258
rect 614 192 617 238
rect 590 142 593 168
rect 622 142 625 278
rect 678 272 681 318
rect 694 312 697 318
rect 718 272 721 518
rect 726 482 729 518
rect 734 482 737 488
rect 734 462 737 478
rect 742 442 745 518
rect 754 478 758 481
rect 750 462 753 468
rect 758 462 761 468
rect 774 452 777 478
rect 774 392 777 448
rect 762 388 766 391
rect 770 368 774 371
rect 726 362 729 368
rect 750 362 753 368
rect 726 302 729 358
rect 782 352 785 538
rect 798 522 801 718
rect 806 702 809 758
rect 830 752 833 778
rect 894 772 897 778
rect 846 752 849 758
rect 854 752 857 758
rect 814 722 817 728
rect 814 692 817 718
rect 830 692 833 698
rect 838 682 841 738
rect 846 702 849 748
rect 862 702 865 768
rect 886 762 889 768
rect 958 762 961 848
rect 966 792 969 848
rect 990 832 993 868
rect 990 792 993 828
rect 978 768 982 771
rect 990 762 993 768
rect 906 758 910 761
rect 890 748 894 751
rect 894 742 897 748
rect 910 712 913 748
rect 918 742 921 748
rect 942 722 945 748
rect 966 732 969 748
rect 874 688 878 691
rect 910 682 913 688
rect 942 682 945 688
rect 822 672 825 678
rect 862 672 865 678
rect 850 668 854 671
rect 890 668 894 671
rect 806 662 809 668
rect 810 658 814 661
rect 850 658 854 661
rect 846 572 849 618
rect 846 562 849 568
rect 862 552 865 668
rect 926 662 929 668
rect 958 662 961 668
rect 902 652 905 658
rect 874 648 878 651
rect 878 582 881 588
rect 902 562 905 648
rect 910 552 913 658
rect 966 632 969 728
rect 980 703 981 707
rect 985 703 986 707
rect 990 703 992 707
rect 998 692 1001 828
rect 1014 742 1017 858
rect 1038 782 1041 868
rect 1062 822 1065 1108
rect 1094 1102 1097 1138
rect 1070 1092 1073 1098
rect 1078 1082 1081 1088
rect 1086 1082 1089 1088
rect 1102 1062 1105 1198
rect 1134 1192 1137 1231
rect 1182 1228 1193 1231
rect 1110 1172 1113 1188
rect 1170 1148 1174 1151
rect 1150 1142 1153 1148
rect 1094 1052 1097 1058
rect 1110 1031 1113 1118
rect 1126 1072 1129 1138
rect 1190 1111 1193 1228
rect 1230 1192 1233 1231
rect 1254 1212 1257 1231
rect 1238 1192 1241 1208
rect 1374 1192 1377 1231
rect 1422 1192 1425 1231
rect 1446 1192 1449 1231
rect 1486 1162 1489 1168
rect 1294 1142 1297 1148
rect 1410 1148 1414 1151
rect 1434 1148 1438 1151
rect 1450 1148 1454 1151
rect 1182 1108 1193 1111
rect 1134 1062 1137 1098
rect 1110 1028 1121 1031
rect 1110 972 1113 1018
rect 1118 962 1121 1028
rect 1134 952 1137 1058
rect 1142 1052 1145 1108
rect 1166 1072 1169 1078
rect 1182 1062 1185 1108
rect 1206 1082 1209 1118
rect 1238 1092 1241 1138
rect 1294 1092 1297 1128
rect 1326 1092 1329 1147
rect 1358 1092 1361 1148
rect 1342 1082 1345 1088
rect 1250 1078 1254 1081
rect 1382 1072 1385 1078
rect 1398 1072 1401 1138
rect 1282 1068 1286 1071
rect 1162 1058 1166 1061
rect 1174 1052 1177 1058
rect 1206 1042 1209 1058
rect 1214 1052 1217 1068
rect 1222 1062 1225 1068
rect 1310 1062 1313 1068
rect 1290 1058 1294 1061
rect 1270 1052 1273 1058
rect 1302 1042 1305 1048
rect 1286 1032 1289 1038
rect 1190 972 1193 1018
rect 1254 972 1257 978
rect 1150 952 1153 958
rect 1086 892 1089 947
rect 1130 938 1134 941
rect 1142 902 1145 938
rect 1150 912 1153 948
rect 1146 888 1150 891
rect 1098 868 1102 871
rect 1070 842 1073 868
rect 1158 862 1161 968
rect 1238 962 1241 968
rect 1166 952 1169 958
rect 1174 952 1177 958
rect 1190 952 1193 958
rect 1218 948 1222 951
rect 1258 948 1262 951
rect 1174 922 1177 938
rect 1166 872 1169 908
rect 1190 872 1193 948
rect 1242 938 1246 941
rect 1254 932 1257 948
rect 1270 942 1273 958
rect 1302 922 1305 947
rect 1242 918 1246 921
rect 1214 892 1217 898
rect 1202 868 1206 871
rect 1082 858 1086 861
rect 1106 858 1110 861
rect 1088 848 1089 851
rect 1098 848 1102 851
rect 1086 842 1089 848
rect 1142 842 1145 858
rect 1166 852 1169 868
rect 1190 862 1193 868
rect 1310 862 1313 1058
rect 1318 1052 1321 1068
rect 1378 1058 1382 1061
rect 1358 1052 1361 1058
rect 1398 982 1401 1068
rect 1418 1058 1422 1061
rect 1422 982 1425 988
rect 1334 952 1337 978
rect 1370 968 1374 971
rect 1366 962 1369 968
rect 1406 952 1409 968
rect 1334 872 1337 948
rect 1378 938 1382 941
rect 1390 932 1393 938
rect 1038 752 1041 758
rect 1038 742 1041 748
rect 1062 742 1065 818
rect 1086 772 1089 778
rect 1074 768 1078 771
rect 1094 762 1097 798
rect 1006 682 1009 688
rect 1038 661 1041 738
rect 1046 672 1049 738
rect 1054 712 1057 728
rect 1054 682 1057 708
rect 1062 672 1065 738
rect 1086 732 1089 748
rect 1094 671 1097 758
rect 1102 742 1105 788
rect 1142 772 1145 778
rect 1166 762 1169 848
rect 1198 842 1201 848
rect 1182 832 1185 838
rect 1150 758 1158 761
rect 1118 752 1121 758
rect 1126 702 1129 758
rect 1138 748 1142 751
rect 1134 722 1137 738
rect 1086 668 1097 671
rect 1122 668 1126 671
rect 1086 662 1089 668
rect 1034 658 1041 661
rect 1050 658 1054 661
rect 1038 652 1041 658
rect 818 548 822 551
rect 806 502 809 548
rect 814 522 817 538
rect 822 522 825 548
rect 870 532 873 538
rect 902 532 905 548
rect 918 542 921 578
rect 942 572 945 628
rect 1038 602 1041 648
rect 1078 642 1081 648
rect 966 592 969 598
rect 926 552 929 558
rect 942 552 945 568
rect 1030 551 1033 588
rect 1062 552 1065 638
rect 934 532 937 538
rect 870 522 873 528
rect 898 518 902 521
rect 830 502 833 508
rect 838 502 841 518
rect 830 492 833 498
rect 794 488 798 491
rect 822 482 825 488
rect 802 448 806 451
rect 814 442 817 468
rect 838 462 841 488
rect 910 472 913 528
rect 980 503 981 507
rect 985 503 986 507
rect 990 503 992 507
rect 882 468 889 471
rect 862 462 865 468
rect 886 462 889 468
rect 842 448 846 451
rect 798 372 801 378
rect 742 342 745 348
rect 758 342 761 348
rect 726 262 729 298
rect 766 282 769 348
rect 790 282 793 368
rect 798 352 801 368
rect 830 332 833 368
rect 846 352 849 358
rect 854 341 857 358
rect 846 338 857 341
rect 814 292 817 318
rect 758 262 761 278
rect 766 272 769 278
rect 642 258 646 261
rect 686 252 689 258
rect 766 251 769 258
rect 762 248 769 251
rect 790 252 793 278
rect 798 272 801 278
rect 654 242 657 248
rect 634 238 638 241
rect 646 212 649 218
rect 642 188 646 191
rect 602 128 606 131
rect 586 68 590 71
rect 462 52 465 58
rect 582 52 585 58
rect 614 52 617 138
rect 630 132 633 168
rect 654 162 657 198
rect 694 182 697 188
rect 662 152 665 158
rect 646 148 654 151
rect 638 142 641 148
rect 630 71 633 128
rect 630 68 638 71
rect 622 62 625 68
rect 646 62 649 148
rect 686 142 689 148
rect 710 142 713 218
rect 722 148 726 151
rect 766 151 769 248
rect 774 202 777 218
rect 766 148 774 151
rect 738 138 742 141
rect 678 132 681 138
rect 706 128 710 131
rect 718 102 721 138
rect 786 128 790 131
rect 750 122 753 128
rect 706 88 710 91
rect 694 62 697 68
rect 674 58 678 61
rect 638 52 641 58
rect 512 48 518 51
rect 666 48 670 51
rect 422 -22 425 48
rect 438 42 441 48
rect 476 3 477 7
rect 481 3 482 7
rect 486 3 488 7
rect 590 -22 593 8
rect 614 -22 617 48
rect 622 42 625 48
rect 690 38 694 41
rect 630 -22 633 8
rect 662 -22 665 18
rect 718 -22 721 98
rect 742 42 745 118
rect 798 92 801 268
rect 810 258 814 261
rect 822 252 825 258
rect 846 252 849 338
rect 862 332 865 458
rect 894 452 897 468
rect 902 462 905 468
rect 910 462 913 468
rect 926 451 929 468
rect 934 462 937 488
rect 966 462 969 468
rect 1006 462 1009 528
rect 1022 482 1025 508
rect 1018 478 1022 481
rect 1002 458 1006 461
rect 958 452 961 458
rect 926 448 934 451
rect 942 442 945 448
rect 886 432 889 438
rect 926 432 929 438
rect 958 432 961 438
rect 898 348 902 351
rect 878 342 881 348
rect 878 292 881 328
rect 894 272 897 328
rect 858 268 862 271
rect 870 262 873 268
rect 842 248 846 251
rect 830 172 833 218
rect 810 148 814 151
rect 846 142 849 248
rect 878 162 881 218
rect 874 148 878 151
rect 810 138 814 141
rect 854 132 857 148
rect 894 142 897 268
rect 910 152 913 388
rect 942 342 945 418
rect 1006 382 1009 458
rect 1046 442 1049 538
rect 1078 532 1081 628
rect 1086 561 1089 658
rect 1094 652 1097 658
rect 1102 632 1105 668
rect 1110 642 1113 658
rect 1126 652 1129 658
rect 1142 642 1145 728
rect 1150 692 1153 758
rect 1190 752 1193 818
rect 1158 662 1161 748
rect 1166 732 1169 748
rect 1198 742 1201 778
rect 1206 752 1209 838
rect 1226 818 1230 821
rect 1294 821 1297 859
rect 1294 818 1305 821
rect 1222 741 1225 768
rect 1230 752 1233 818
rect 1246 762 1249 768
rect 1248 758 1249 762
rect 1222 738 1230 741
rect 1182 732 1185 738
rect 1174 712 1177 718
rect 1166 682 1169 708
rect 1150 652 1153 658
rect 1158 652 1161 658
rect 1166 642 1169 678
rect 1190 661 1193 738
rect 1230 732 1233 738
rect 1222 672 1225 718
rect 1246 682 1249 688
rect 1254 672 1257 758
rect 1266 748 1270 751
rect 1262 732 1265 738
rect 1270 681 1273 748
rect 1294 692 1297 798
rect 1302 792 1305 818
rect 1302 752 1305 768
rect 1318 762 1321 768
rect 1326 742 1329 838
rect 1350 802 1353 859
rect 1366 752 1369 758
rect 1302 682 1305 728
rect 1342 722 1345 738
rect 1350 722 1353 748
rect 1374 732 1377 928
rect 1382 772 1385 778
rect 1398 752 1401 948
rect 1430 942 1433 948
rect 1438 932 1441 958
rect 1446 952 1449 1148
rect 1474 1088 1478 1091
rect 1446 932 1449 948
rect 1430 892 1433 928
rect 1418 838 1422 841
rect 1430 772 1433 818
rect 1446 812 1449 858
rect 1454 842 1457 858
rect 1334 712 1337 718
rect 1334 702 1337 708
rect 1262 678 1273 681
rect 1262 672 1265 678
rect 1278 671 1281 678
rect 1274 668 1281 671
rect 1302 672 1305 678
rect 1322 668 1326 671
rect 1230 662 1233 668
rect 1186 658 1193 661
rect 1202 658 1206 661
rect 1174 652 1177 658
rect 1246 652 1249 668
rect 1334 662 1337 678
rect 1358 672 1361 688
rect 1366 672 1369 708
rect 1374 662 1377 718
rect 1382 682 1385 748
rect 1402 728 1406 731
rect 1414 721 1417 758
rect 1426 748 1430 751
rect 1438 742 1441 748
rect 1406 718 1417 721
rect 1390 682 1393 688
rect 1406 682 1409 718
rect 1398 672 1401 678
rect 1406 662 1409 668
rect 1258 658 1262 661
rect 1282 658 1286 661
rect 1330 658 1334 661
rect 1378 658 1382 661
rect 1186 648 1190 651
rect 1298 648 1302 651
rect 1338 648 1344 651
rect 1198 622 1201 628
rect 1102 592 1105 608
rect 1086 558 1097 561
rect 1086 522 1089 548
rect 1030 412 1033 418
rect 1054 362 1057 378
rect 1040 358 1046 361
rect 986 348 990 351
rect 1010 348 1014 351
rect 1022 342 1025 358
rect 1062 352 1065 378
rect 1070 372 1073 518
rect 1034 348 1038 351
rect 994 338 998 341
rect 918 262 921 338
rect 934 292 937 328
rect 942 272 945 338
rect 1022 332 1025 338
rect 1054 332 1057 338
rect 980 303 981 307
rect 985 303 986 307
rect 990 303 992 307
rect 942 262 945 268
rect 942 152 945 178
rect 966 162 969 278
rect 982 262 985 288
rect 1078 272 1081 468
rect 1086 442 1089 458
rect 1094 392 1097 558
rect 1118 532 1121 558
rect 1126 472 1129 598
rect 1190 582 1193 588
rect 1134 572 1137 578
rect 1134 492 1137 548
rect 1142 542 1145 558
rect 1190 552 1193 568
rect 1154 548 1158 551
rect 1142 462 1145 518
rect 1206 482 1209 638
rect 1214 562 1217 588
rect 1246 582 1249 648
rect 1254 572 1257 578
rect 1294 572 1297 638
rect 1302 592 1305 618
rect 1334 592 1337 638
rect 1230 541 1233 568
rect 1238 552 1241 558
rect 1302 552 1305 558
rect 1358 552 1361 658
rect 1394 648 1398 651
rect 1398 572 1401 578
rect 1406 552 1409 658
rect 1414 652 1417 658
rect 1422 641 1425 738
rect 1446 682 1449 778
rect 1430 652 1433 678
rect 1454 662 1457 768
rect 1422 638 1433 641
rect 1422 572 1425 598
rect 1246 542 1249 548
rect 1254 542 1257 548
rect 1278 542 1281 548
rect 1230 538 1238 541
rect 1274 538 1278 541
rect 1182 462 1185 468
rect 1142 421 1145 458
rect 1142 418 1153 421
rect 1110 362 1113 368
rect 1094 352 1097 358
rect 1102 352 1105 358
rect 1142 351 1145 358
rect 1126 342 1129 348
rect 1078 262 1081 268
rect 1026 258 1030 261
rect 1106 259 1110 261
rect 1106 258 1113 259
rect 1142 242 1145 278
rect 1050 238 1054 241
rect 1014 162 1017 218
rect 1006 152 1009 158
rect 1014 142 1017 148
rect 978 138 982 141
rect 1038 141 1041 218
rect 1110 152 1113 158
rect 1058 148 1062 151
rect 1082 148 1086 151
rect 1102 142 1105 148
rect 1038 138 1046 141
rect 958 132 961 138
rect 938 128 942 131
rect 1022 122 1025 128
rect 866 118 870 121
rect 806 82 809 118
rect 782 62 785 68
rect 814 62 817 78
rect 838 62 841 98
rect 878 62 881 118
rect 926 82 929 118
rect 950 102 953 118
rect 980 103 981 107
rect 985 103 986 107
rect 990 103 992 107
rect 1038 92 1041 128
rect 934 82 937 88
rect 902 62 905 68
rect 754 58 758 61
rect 1042 58 1046 61
rect 966 42 969 58
rect 1062 42 1065 128
rect 1070 82 1073 108
rect 1070 63 1073 68
rect 1086 62 1089 138
rect 1142 132 1145 238
rect 1150 152 1153 418
rect 1158 362 1161 418
rect 1206 392 1209 478
rect 1214 462 1217 468
rect 1246 462 1249 538
rect 1302 512 1305 548
rect 1314 538 1318 541
rect 1322 528 1326 531
rect 1266 488 1270 491
rect 1302 482 1305 488
rect 1290 468 1294 471
rect 1318 471 1321 518
rect 1358 512 1361 548
rect 1374 541 1377 548
rect 1366 538 1377 541
rect 1318 468 1329 471
rect 1278 462 1281 468
rect 1266 458 1270 461
rect 1314 458 1318 461
rect 1206 382 1209 388
rect 1214 352 1217 388
rect 1278 362 1281 458
rect 1326 452 1329 468
rect 1334 392 1337 498
rect 1342 462 1345 508
rect 1366 481 1369 538
rect 1374 522 1377 528
rect 1362 478 1369 481
rect 1354 468 1358 471
rect 1382 462 1385 548
rect 1406 542 1409 548
rect 1394 468 1398 471
rect 1406 462 1409 488
rect 1414 452 1417 518
rect 1422 502 1425 548
rect 1430 532 1433 638
rect 1438 542 1441 618
rect 1462 592 1465 1038
rect 1486 992 1489 998
rect 1486 862 1489 868
rect 1486 792 1489 798
rect 1446 582 1449 588
rect 1454 542 1457 548
rect 1454 492 1457 528
rect 1470 482 1473 718
rect 1478 572 1481 738
rect 1486 692 1489 698
rect 1422 462 1425 468
rect 1438 458 1446 461
rect 1402 448 1406 451
rect 1342 372 1345 418
rect 1222 342 1225 358
rect 1282 348 1286 351
rect 1338 348 1342 351
rect 1254 342 1257 348
rect 1238 322 1241 328
rect 1190 272 1193 278
rect 1158 262 1161 268
rect 1230 262 1233 318
rect 1286 292 1289 328
rect 1318 292 1321 348
rect 1350 342 1353 358
rect 1366 352 1369 418
rect 1398 392 1401 438
rect 1430 382 1433 388
rect 1374 352 1377 358
rect 1438 352 1441 458
rect 1486 362 1489 368
rect 1334 292 1337 318
rect 1358 292 1361 318
rect 1270 282 1273 288
rect 1350 282 1353 288
rect 1298 278 1302 281
rect 1366 272 1369 338
rect 1406 332 1409 338
rect 1414 332 1417 348
rect 1394 328 1398 331
rect 1438 322 1441 348
rect 1446 292 1449 328
rect 1302 262 1305 268
rect 1310 262 1313 268
rect 1274 258 1278 261
rect 1330 258 1334 261
rect 1174 142 1177 258
rect 1206 152 1209 168
rect 1214 152 1217 158
rect 1230 142 1233 148
rect 1246 132 1249 168
rect 1102 62 1105 128
rect 1190 101 1193 118
rect 1190 98 1201 101
rect 1198 62 1201 98
rect 1246 62 1249 128
rect 1270 72 1273 258
rect 1290 148 1294 151
rect 1302 92 1305 148
rect 1374 142 1377 147
rect 1382 142 1385 268
rect 1390 262 1393 288
rect 1454 262 1457 278
rect 1442 148 1446 151
rect 1434 118 1438 121
rect 1318 72 1321 118
rect 1454 92 1457 248
rect 1462 192 1465 318
rect 1486 262 1489 268
rect 1446 72 1449 78
rect 1462 62 1465 118
rect 1070 58 1073 59
rect 1130 58 1134 61
rect 1154 58 1158 61
rect 1178 58 1182 61
rect 1218 58 1222 61
rect 1378 58 1382 61
rect 1402 58 1406 61
rect 1426 58 1430 61
rect 1486 52 1489 158
rect 1002 38 1006 41
rect 798 -22 801 18
rect 822 -22 825 18
rect 886 -22 889 8
rect 918 -22 921 8
rect 958 -22 961 18
rect 982 -22 985 18
rect 1022 -22 1025 8
rect 1038 -22 1041 8
rect 1118 -22 1121 18
rect 1142 -22 1145 18
rect 1214 -22 1217 18
rect 1262 -22 1265 18
rect 1342 -22 1345 18
rect 1390 -22 1393 18
rect 1414 -22 1417 18
rect 1438 -22 1441 18
<< m3contact >>
rect 166 1208 170 1212
rect 472 1203 476 1207
rect 477 1203 481 1207
rect 482 1203 486 1207
rect 614 1208 618 1212
rect 198 1168 202 1172
rect 214 1168 218 1172
rect 318 1168 322 1172
rect 70 1158 74 1162
rect 142 1158 146 1162
rect 174 1148 178 1152
rect 6 1128 10 1132
rect 126 1128 130 1132
rect 174 1128 178 1132
rect 190 1128 194 1132
rect 62 1068 66 1072
rect 166 1108 170 1112
rect 406 1158 410 1162
rect 422 1158 426 1162
rect 638 1158 642 1162
rect 654 1158 658 1162
rect 662 1158 666 1162
rect 734 1158 738 1162
rect 390 1148 394 1152
rect 414 1148 418 1152
rect 382 1138 386 1142
rect 366 1128 370 1132
rect 286 1108 290 1112
rect 334 1108 338 1112
rect 374 1108 378 1112
rect 406 1118 410 1122
rect 438 1148 442 1152
rect 526 1148 530 1152
rect 454 1138 458 1142
rect 446 1128 450 1132
rect 430 1108 434 1112
rect 286 1078 290 1082
rect 398 1078 402 1082
rect 126 1068 130 1072
rect 198 1068 202 1072
rect 374 1068 378 1072
rect 6 1058 10 1062
rect 86 1058 90 1062
rect 142 1058 146 1062
rect 6 988 10 992
rect 22 968 26 972
rect 142 968 146 972
rect 30 958 34 962
rect 134 948 138 952
rect 46 888 50 892
rect 118 918 122 922
rect 142 918 146 922
rect 190 968 194 972
rect 182 938 186 942
rect 158 898 162 902
rect 126 878 130 882
rect 62 868 66 872
rect 6 858 10 862
rect 6 758 10 762
rect 214 958 218 962
rect 254 1048 258 1052
rect 286 1048 290 1052
rect 334 1038 338 1042
rect 518 1118 522 1122
rect 462 1078 466 1082
rect 558 1128 562 1132
rect 550 1118 554 1122
rect 542 1108 546 1112
rect 582 1118 586 1122
rect 598 1118 602 1122
rect 630 1108 634 1112
rect 526 1078 530 1082
rect 470 1068 474 1072
rect 510 1068 514 1072
rect 558 1068 562 1072
rect 582 1068 586 1072
rect 614 1068 618 1072
rect 414 1058 418 1062
rect 430 1058 434 1062
rect 454 1058 458 1062
rect 590 1058 594 1062
rect 622 1058 626 1062
rect 246 968 250 972
rect 398 968 402 972
rect 262 958 266 962
rect 318 958 322 962
rect 438 1048 442 1052
rect 430 968 434 972
rect 294 948 298 952
rect 318 948 322 952
rect 326 948 330 952
rect 358 948 362 952
rect 326 938 330 942
rect 358 928 362 932
rect 406 928 410 932
rect 270 918 274 922
rect 302 918 306 922
rect 246 908 250 912
rect 446 1038 450 1042
rect 438 958 442 962
rect 472 1003 476 1007
rect 477 1003 481 1007
rect 482 1003 486 1007
rect 454 948 458 952
rect 566 1048 570 1052
rect 590 1048 594 1052
rect 614 1038 618 1042
rect 590 968 594 972
rect 574 958 578 962
rect 510 948 514 952
rect 550 948 554 952
rect 430 938 434 942
rect 414 918 418 922
rect 334 908 338 912
rect 286 888 290 892
rect 230 868 234 872
rect 182 858 186 862
rect 246 858 250 862
rect 94 838 98 842
rect 134 828 138 832
rect 126 768 130 772
rect 214 848 218 852
rect 190 828 194 832
rect 350 878 354 882
rect 462 888 466 892
rect 334 858 338 862
rect 430 858 434 862
rect 446 858 450 862
rect 470 868 474 872
rect 486 858 490 862
rect 526 938 530 942
rect 534 918 538 922
rect 534 888 538 892
rect 510 878 514 882
rect 558 938 562 942
rect 654 1058 658 1062
rect 638 1048 642 1052
rect 646 1048 650 1052
rect 630 958 634 962
rect 646 958 650 962
rect 622 948 626 952
rect 630 948 634 952
rect 574 928 578 932
rect 582 918 586 922
rect 566 888 570 892
rect 622 928 626 932
rect 622 888 626 892
rect 598 878 602 882
rect 646 878 650 882
rect 574 868 578 872
rect 542 858 546 862
rect 278 848 282 852
rect 454 848 458 852
rect 494 848 498 852
rect 222 818 226 822
rect 158 758 162 762
rect 166 758 170 762
rect 310 838 314 842
rect 342 838 346 842
rect 438 838 442 842
rect 438 828 442 832
rect 478 828 482 832
rect 472 803 476 807
rect 477 803 481 807
rect 482 803 486 807
rect 534 838 538 842
rect 518 828 522 832
rect 358 778 362 782
rect 510 778 514 782
rect 246 768 250 772
rect 70 748 74 752
rect 134 748 138 752
rect 62 738 66 742
rect 38 728 42 732
rect 54 728 58 732
rect 94 728 98 732
rect 38 668 42 672
rect 6 658 10 662
rect 118 738 122 742
rect 254 758 258 762
rect 310 758 314 762
rect 238 738 242 742
rect 302 748 306 752
rect 278 738 282 742
rect 158 728 162 732
rect 206 728 210 732
rect 230 728 234 732
rect 246 728 250 732
rect 254 728 258 732
rect 286 728 290 732
rect 294 728 298 732
rect 310 728 314 732
rect 102 718 106 722
rect 126 718 130 722
rect 70 688 74 692
rect 174 698 178 702
rect 206 698 210 702
rect 126 678 130 682
rect 190 678 194 682
rect 222 678 226 682
rect 142 668 146 672
rect 94 648 98 652
rect 6 588 10 592
rect 62 588 66 592
rect 86 588 90 592
rect 206 658 210 662
rect 254 718 258 722
rect 254 688 258 692
rect 270 688 274 692
rect 254 658 258 662
rect 158 648 162 652
rect 190 588 194 592
rect 30 558 34 562
rect 158 558 162 562
rect 54 548 58 552
rect 94 548 98 552
rect 126 548 130 552
rect 6 528 10 532
rect 22 528 26 532
rect 46 528 50 532
rect 62 488 66 492
rect 102 488 106 492
rect 86 478 90 482
rect 70 468 74 472
rect 102 468 106 472
rect 118 468 122 472
rect 6 358 10 362
rect 278 668 282 672
rect 318 718 322 722
rect 326 718 330 722
rect 326 668 330 672
rect 334 668 338 672
rect 390 768 394 772
rect 406 768 410 772
rect 462 758 466 762
rect 422 748 426 752
rect 374 738 378 742
rect 366 728 370 732
rect 398 738 402 742
rect 430 738 434 742
rect 462 738 466 742
rect 398 728 402 732
rect 382 718 386 722
rect 518 748 522 752
rect 502 738 506 742
rect 454 728 458 732
rect 582 858 586 862
rect 566 848 570 852
rect 582 848 586 852
rect 590 848 594 852
rect 574 778 578 782
rect 566 748 570 752
rect 550 738 554 742
rect 542 728 546 732
rect 486 718 490 722
rect 518 718 522 722
rect 542 698 546 702
rect 550 688 554 692
rect 430 678 434 682
rect 542 678 546 682
rect 374 668 378 672
rect 398 668 402 672
rect 414 668 418 672
rect 358 658 362 662
rect 406 658 410 662
rect 350 648 354 652
rect 382 648 386 652
rect 430 648 434 652
rect 270 638 274 642
rect 334 638 338 642
rect 390 618 394 622
rect 310 588 314 592
rect 342 578 346 582
rect 238 558 242 562
rect 214 548 218 552
rect 398 588 402 592
rect 350 548 354 552
rect 366 548 370 552
rect 174 538 178 542
rect 254 528 258 532
rect 230 518 234 522
rect 270 518 274 522
rect 302 518 306 522
rect 182 498 186 502
rect 174 478 178 482
rect 158 468 162 472
rect 126 448 130 452
rect 134 378 138 382
rect 94 358 98 362
rect 62 338 66 342
rect 126 338 130 342
rect 6 298 10 302
rect 70 268 74 272
rect 102 258 106 262
rect 166 448 170 452
rect 198 468 202 472
rect 206 468 210 472
rect 206 448 210 452
rect 190 438 194 442
rect 254 498 258 502
rect 246 478 250 482
rect 286 478 290 482
rect 238 378 242 382
rect 230 368 234 372
rect 142 348 146 352
rect 198 348 202 352
rect 222 348 226 352
rect 174 338 178 342
rect 174 318 178 322
rect 118 248 122 252
rect 110 188 114 192
rect 110 168 114 172
rect 86 148 90 152
rect 62 128 66 132
rect 14 118 18 122
rect 22 118 26 122
rect 94 108 98 112
rect 70 88 74 92
rect 30 78 34 82
rect 86 78 90 82
rect 38 68 42 72
rect 102 78 106 82
rect 6 58 10 62
rect 54 58 58 62
rect 78 58 82 62
rect 174 258 178 262
rect 214 338 218 342
rect 206 288 210 292
rect 198 278 202 282
rect 310 498 314 502
rect 254 458 258 462
rect 366 508 370 512
rect 550 658 554 662
rect 486 648 490 652
rect 470 638 474 642
rect 534 638 538 642
rect 558 638 562 642
rect 414 558 418 562
rect 574 648 578 652
rect 472 603 476 607
rect 477 603 481 607
rect 482 603 486 607
rect 542 578 546 582
rect 422 548 426 552
rect 438 548 442 552
rect 470 548 474 552
rect 550 548 554 552
rect 406 538 410 542
rect 542 538 546 542
rect 398 528 402 532
rect 494 528 498 532
rect 422 508 426 512
rect 342 468 346 472
rect 334 458 338 462
rect 278 448 282 452
rect 262 438 266 442
rect 254 358 258 362
rect 278 358 282 362
rect 286 348 290 352
rect 286 328 290 332
rect 246 298 250 302
rect 270 288 274 292
rect 206 258 210 262
rect 190 248 194 252
rect 166 188 170 192
rect 134 168 138 172
rect 246 238 250 242
rect 206 178 210 182
rect 134 158 138 162
rect 166 158 170 162
rect 166 118 170 122
rect 270 218 274 222
rect 278 188 282 192
rect 254 168 258 172
rect 198 158 202 162
rect 222 148 226 152
rect 206 138 210 142
rect 182 108 186 112
rect 182 98 186 102
rect 118 88 122 92
rect 158 88 162 92
rect 158 78 162 82
rect 262 158 266 162
rect 238 138 242 142
rect 214 128 218 132
rect 238 108 242 112
rect 238 98 242 102
rect 222 88 226 92
rect 206 78 210 82
rect 126 68 130 72
rect 182 58 186 62
rect 230 58 234 62
rect 286 178 290 182
rect 342 438 346 442
rect 358 388 362 392
rect 342 378 346 382
rect 326 358 330 362
rect 446 458 450 462
rect 430 448 434 452
rect 678 1128 682 1132
rect 854 1148 858 1152
rect 790 1138 794 1142
rect 750 1108 754 1112
rect 782 1108 786 1112
rect 678 1088 682 1092
rect 686 1088 690 1092
rect 742 1088 746 1092
rect 670 1078 674 1082
rect 670 1058 674 1062
rect 726 1048 730 1052
rect 798 1058 802 1062
rect 686 998 690 1002
rect 678 948 682 952
rect 678 938 682 942
rect 646 868 650 872
rect 654 868 658 872
rect 606 858 610 862
rect 630 858 634 862
rect 654 848 658 852
rect 622 788 626 792
rect 598 768 602 772
rect 750 958 754 962
rect 710 948 714 952
rect 814 998 818 1002
rect 702 928 706 932
rect 718 898 722 902
rect 750 888 754 892
rect 822 938 826 942
rect 774 878 778 882
rect 782 878 786 882
rect 694 868 698 872
rect 718 868 722 872
rect 742 858 746 862
rect 686 838 690 842
rect 718 808 722 812
rect 822 848 826 852
rect 678 778 682 782
rect 774 778 778 782
rect 790 778 794 782
rect 694 758 698 762
rect 662 748 666 752
rect 590 698 594 702
rect 710 718 714 722
rect 726 718 730 722
rect 726 708 730 712
rect 766 698 770 702
rect 606 688 610 692
rect 598 648 602 652
rect 702 678 706 682
rect 622 668 626 672
rect 646 668 650 672
rect 846 998 850 1002
rect 870 1208 874 1212
rect 886 1208 890 1212
rect 894 1208 898 1212
rect 910 1208 914 1212
rect 918 1208 922 1212
rect 934 1208 938 1212
rect 998 1208 1002 1212
rect 1038 1208 1042 1212
rect 1054 1208 1058 1212
rect 1062 1208 1066 1212
rect 1078 1208 1082 1212
rect 1102 1198 1106 1202
rect 1118 1198 1122 1202
rect 870 1148 874 1152
rect 894 1148 898 1152
rect 878 1108 882 1112
rect 926 1088 930 1092
rect 974 1118 978 1122
rect 1014 1118 1018 1122
rect 976 1103 980 1107
rect 981 1103 985 1107
rect 986 1103 990 1107
rect 950 1088 954 1092
rect 926 1068 930 1072
rect 1078 1138 1082 1142
rect 1094 1138 1098 1142
rect 1046 1108 1050 1112
rect 1062 1108 1066 1112
rect 1086 1108 1090 1112
rect 1022 1098 1026 1102
rect 1054 1068 1058 1072
rect 990 1058 994 1062
rect 966 1048 970 1052
rect 998 1008 1002 1012
rect 902 968 906 972
rect 910 958 914 962
rect 942 948 946 952
rect 854 938 858 942
rect 862 938 866 942
rect 894 938 898 942
rect 918 938 922 942
rect 974 928 978 932
rect 966 918 970 922
rect 838 888 842 892
rect 878 888 882 892
rect 1030 908 1034 912
rect 976 903 980 907
rect 981 903 985 907
rect 986 903 990 907
rect 862 878 866 882
rect 950 878 954 882
rect 1054 908 1058 912
rect 950 868 954 872
rect 942 858 946 862
rect 870 828 874 832
rect 934 838 938 842
rect 878 808 882 812
rect 958 848 962 852
rect 982 848 986 852
rect 942 818 946 822
rect 830 788 834 792
rect 830 778 834 782
rect 814 768 818 772
rect 798 758 802 762
rect 790 728 794 732
rect 702 658 706 662
rect 630 638 634 642
rect 582 568 586 572
rect 774 648 778 652
rect 790 668 794 672
rect 782 618 786 622
rect 782 608 786 612
rect 646 548 650 552
rect 694 548 698 552
rect 710 548 714 552
rect 606 538 610 542
rect 638 538 642 542
rect 686 538 690 542
rect 702 538 706 542
rect 654 528 658 532
rect 630 518 634 522
rect 646 498 650 502
rect 614 478 618 482
rect 630 478 634 482
rect 654 478 658 482
rect 670 478 674 482
rect 646 468 650 472
rect 566 448 570 452
rect 638 448 642 452
rect 574 438 578 442
rect 598 438 602 442
rect 534 418 538 422
rect 472 403 476 407
rect 477 403 481 407
rect 482 403 486 407
rect 526 388 530 392
rect 550 388 554 392
rect 406 368 410 372
rect 374 358 378 362
rect 518 358 522 362
rect 342 348 346 352
rect 398 348 402 352
rect 302 338 306 342
rect 366 338 370 342
rect 438 338 442 342
rect 326 328 330 332
rect 310 308 314 312
rect 318 298 322 302
rect 462 348 466 352
rect 534 348 538 352
rect 438 328 442 332
rect 454 328 458 332
rect 422 318 426 322
rect 430 318 434 322
rect 374 308 378 312
rect 310 268 314 272
rect 358 268 362 272
rect 326 238 330 242
rect 310 228 314 232
rect 326 188 330 192
rect 302 168 306 172
rect 286 148 290 152
rect 310 158 314 162
rect 350 148 354 152
rect 318 138 322 142
rect 390 288 394 292
rect 414 278 418 282
rect 382 268 386 272
rect 422 268 426 272
rect 398 248 402 252
rect 374 148 378 152
rect 366 138 370 142
rect 366 128 370 132
rect 270 118 274 122
rect 366 108 370 112
rect 350 98 354 102
rect 294 88 298 92
rect 398 158 402 162
rect 382 88 386 92
rect 358 78 362 82
rect 286 68 290 72
rect 294 58 298 62
rect 326 58 330 62
rect 158 48 162 52
rect 190 48 194 52
rect 254 48 258 52
rect 310 38 314 42
rect 438 278 442 282
rect 462 308 466 312
rect 462 298 466 302
rect 582 378 586 382
rect 582 348 586 352
rect 558 338 562 342
rect 518 328 522 332
rect 574 328 578 332
rect 518 298 522 302
rect 510 278 514 282
rect 542 278 546 282
rect 446 268 450 272
rect 542 268 546 272
rect 574 268 578 272
rect 446 258 450 262
rect 502 258 506 262
rect 526 258 530 262
rect 566 258 570 262
rect 630 378 634 382
rect 614 368 618 372
rect 606 348 610 352
rect 598 328 602 332
rect 598 318 602 322
rect 606 318 610 322
rect 598 278 602 282
rect 590 268 594 272
rect 758 538 762 542
rect 742 528 746 532
rect 766 528 770 532
rect 718 518 722 522
rect 726 518 730 522
rect 774 518 778 522
rect 694 498 698 502
rect 710 478 714 482
rect 686 458 690 462
rect 670 378 674 382
rect 638 338 642 342
rect 694 348 698 352
rect 662 328 666 332
rect 678 328 682 332
rect 686 328 690 332
rect 710 328 714 332
rect 678 318 682 322
rect 654 278 658 282
rect 478 238 482 242
rect 494 238 498 242
rect 478 228 482 232
rect 486 228 490 232
rect 486 218 490 222
rect 472 203 476 207
rect 477 203 481 207
rect 482 203 486 207
rect 422 168 426 172
rect 414 138 418 142
rect 406 108 410 112
rect 430 158 434 162
rect 454 158 458 162
rect 478 158 482 162
rect 470 138 474 142
rect 454 128 458 132
rect 430 108 434 112
rect 614 258 618 262
rect 518 248 522 252
rect 582 248 586 252
rect 598 248 602 252
rect 558 238 562 242
rect 574 238 578 242
rect 550 228 554 232
rect 518 188 522 192
rect 526 178 530 182
rect 550 178 554 182
rect 542 158 546 162
rect 558 168 562 172
rect 574 168 578 172
rect 526 128 530 132
rect 518 118 522 122
rect 494 108 498 112
rect 510 108 514 112
rect 438 98 442 102
rect 478 98 482 102
rect 470 88 474 92
rect 422 78 426 82
rect 438 68 442 72
rect 422 58 426 62
rect 486 68 490 72
rect 558 118 562 122
rect 566 98 570 102
rect 534 88 538 92
rect 550 78 554 82
rect 590 188 594 192
rect 614 238 618 242
rect 590 168 594 172
rect 606 168 610 172
rect 694 308 698 312
rect 734 488 738 492
rect 734 458 738 462
rect 758 478 762 482
rect 750 468 754 472
rect 758 468 762 472
rect 774 448 778 452
rect 742 438 746 442
rect 766 388 770 392
rect 774 388 778 392
rect 726 368 730 372
rect 750 368 754 372
rect 774 368 778 372
rect 894 768 898 772
rect 854 758 858 762
rect 846 748 850 752
rect 814 728 818 732
rect 814 718 818 722
rect 806 698 810 702
rect 830 698 834 702
rect 1014 858 1018 862
rect 990 828 994 832
rect 998 828 1002 832
rect 990 788 994 792
rect 982 768 986 772
rect 990 768 994 772
rect 886 758 890 762
rect 910 758 914 762
rect 886 748 890 752
rect 910 748 914 752
rect 894 738 898 742
rect 918 738 922 742
rect 966 728 970 732
rect 942 718 946 722
rect 910 708 914 712
rect 846 698 850 702
rect 862 698 866 702
rect 870 688 874 692
rect 910 688 914 692
rect 942 688 946 692
rect 838 678 842 682
rect 862 678 866 682
rect 822 668 826 672
rect 846 668 850 672
rect 894 668 898 672
rect 926 668 930 672
rect 958 668 962 672
rect 814 658 818 662
rect 854 658 858 662
rect 846 618 850 622
rect 846 568 850 572
rect 902 658 906 662
rect 870 648 874 652
rect 878 588 882 592
rect 902 558 906 562
rect 976 703 980 707
rect 981 703 985 707
rect 986 703 990 707
rect 1070 1098 1074 1102
rect 1094 1098 1098 1102
rect 1078 1088 1082 1092
rect 1086 1088 1090 1092
rect 1110 1188 1114 1192
rect 1134 1188 1138 1192
rect 1174 1148 1178 1152
rect 1150 1138 1154 1142
rect 1094 1048 1098 1052
rect 1142 1108 1146 1112
rect 1238 1208 1242 1212
rect 1254 1208 1258 1212
rect 1486 1158 1490 1162
rect 1414 1148 1418 1152
rect 1438 1148 1442 1152
rect 1446 1148 1450 1152
rect 1238 1138 1242 1142
rect 1294 1138 1298 1142
rect 1134 1098 1138 1102
rect 1126 1068 1130 1072
rect 1134 1058 1138 1062
rect 1110 968 1114 972
rect 1166 1078 1170 1082
rect 1166 1068 1170 1072
rect 1398 1138 1402 1142
rect 1294 1088 1298 1092
rect 1342 1088 1346 1092
rect 1358 1088 1362 1092
rect 1206 1078 1210 1082
rect 1246 1078 1250 1082
rect 1222 1068 1226 1072
rect 1286 1068 1290 1072
rect 1310 1068 1314 1072
rect 1382 1068 1386 1072
rect 1166 1058 1170 1062
rect 1174 1048 1178 1052
rect 1294 1058 1298 1062
rect 1214 1048 1218 1052
rect 1270 1048 1274 1052
rect 1206 1038 1210 1042
rect 1302 1038 1306 1042
rect 1286 1028 1290 1032
rect 1254 978 1258 982
rect 1158 968 1162 972
rect 1190 968 1194 972
rect 1238 968 1242 972
rect 1150 948 1154 952
rect 1134 938 1138 942
rect 1150 908 1154 912
rect 1142 898 1146 902
rect 1086 888 1090 892
rect 1150 888 1154 892
rect 1070 868 1074 872
rect 1094 868 1098 872
rect 1174 958 1178 962
rect 1190 958 1194 962
rect 1166 948 1170 952
rect 1214 948 1218 952
rect 1262 948 1266 952
rect 1174 918 1178 922
rect 1166 908 1170 912
rect 1238 938 1242 942
rect 1270 938 1274 942
rect 1254 928 1258 932
rect 1246 918 1250 922
rect 1302 918 1306 922
rect 1214 898 1218 902
rect 1190 868 1194 872
rect 1198 868 1202 872
rect 1086 858 1090 862
rect 1102 858 1106 862
rect 1102 848 1106 852
rect 1374 1058 1378 1062
rect 1318 1048 1322 1052
rect 1358 1048 1362 1052
rect 1414 1058 1418 1062
rect 1422 988 1426 992
rect 1334 978 1338 982
rect 1398 978 1402 982
rect 1374 968 1378 972
rect 1406 968 1410 972
rect 1366 958 1370 962
rect 1438 958 1442 962
rect 1398 948 1402 952
rect 1430 948 1434 952
rect 1382 938 1386 942
rect 1390 928 1394 932
rect 1166 848 1170 852
rect 1070 838 1074 842
rect 1086 838 1090 842
rect 1142 838 1146 842
rect 1062 818 1066 822
rect 1038 778 1042 782
rect 1038 758 1042 762
rect 1094 798 1098 802
rect 1086 778 1090 782
rect 1070 768 1074 772
rect 1102 788 1106 792
rect 1014 738 1018 742
rect 1038 738 1042 742
rect 1006 688 1010 692
rect 1054 708 1058 712
rect 1054 678 1058 682
rect 1086 728 1090 732
rect 1142 778 1146 782
rect 1198 838 1202 842
rect 1206 838 1210 842
rect 1182 828 1186 832
rect 1118 758 1122 762
rect 1166 758 1170 762
rect 1134 748 1138 752
rect 1142 728 1146 732
rect 1134 718 1138 722
rect 1126 698 1130 702
rect 1118 668 1122 672
rect 1054 658 1058 662
rect 1094 658 1098 662
rect 1078 648 1082 652
rect 942 628 946 632
rect 966 628 970 632
rect 918 578 922 582
rect 822 548 826 552
rect 862 548 866 552
rect 902 548 906 552
rect 798 518 802 522
rect 1062 638 1066 642
rect 966 598 970 602
rect 1038 598 1042 602
rect 1030 588 1034 592
rect 942 568 946 572
rect 926 558 930 562
rect 1078 628 1082 632
rect 910 528 914 532
rect 934 528 938 532
rect 1006 528 1010 532
rect 814 518 818 522
rect 822 518 826 522
rect 870 518 874 522
rect 902 518 906 522
rect 830 508 834 512
rect 806 498 810 502
rect 830 498 834 502
rect 838 498 842 502
rect 790 488 794 492
rect 822 488 826 492
rect 838 488 842 492
rect 798 448 802 452
rect 976 503 980 507
rect 981 503 985 507
rect 986 503 990 507
rect 934 488 938 492
rect 878 468 882 472
rect 902 468 906 472
rect 862 458 866 462
rect 838 448 842 452
rect 814 438 818 442
rect 798 378 802 382
rect 790 368 794 372
rect 798 368 802 372
rect 830 368 834 372
rect 742 348 746 352
rect 766 348 770 352
rect 782 348 786 352
rect 758 338 762 342
rect 726 298 730 302
rect 718 268 722 272
rect 846 358 850 362
rect 814 288 818 292
rect 758 278 762 282
rect 766 278 770 282
rect 798 278 802 282
rect 638 258 642 262
rect 758 258 762 262
rect 686 248 690 252
rect 790 248 794 252
rect 630 238 634 242
rect 654 238 658 242
rect 646 208 650 212
rect 654 198 658 202
rect 638 188 642 192
rect 630 168 634 172
rect 614 138 618 142
rect 622 138 626 142
rect 598 128 602 132
rect 582 68 586 72
rect 534 58 538 62
rect 694 188 698 192
rect 662 158 666 162
rect 638 148 642 152
rect 654 148 658 152
rect 718 148 722 152
rect 774 198 778 202
rect 678 138 682 142
rect 686 138 690 142
rect 710 138 714 142
rect 734 138 738 142
rect 702 128 706 132
rect 782 128 786 132
rect 750 118 754 122
rect 718 98 722 102
rect 710 88 714 92
rect 694 68 698 72
rect 622 58 626 62
rect 670 58 674 62
rect 438 48 442 52
rect 462 48 466 52
rect 518 48 522 52
rect 582 48 586 52
rect 638 48 642 52
rect 662 48 666 52
rect 590 8 594 12
rect 472 3 476 7
rect 477 3 481 7
rect 482 3 486 7
rect 622 38 626 42
rect 694 38 698 42
rect 630 8 634 12
rect 814 258 818 262
rect 822 258 826 262
rect 910 458 914 462
rect 894 448 898 452
rect 966 468 970 472
rect 1022 508 1026 512
rect 1014 478 1018 482
rect 998 458 1002 462
rect 934 448 938 452
rect 958 448 962 452
rect 942 438 946 442
rect 886 428 890 432
rect 926 428 930 432
rect 958 428 962 432
rect 942 418 946 422
rect 910 388 914 392
rect 894 348 898 352
rect 878 338 882 342
rect 862 328 866 332
rect 878 328 882 332
rect 854 268 858 272
rect 894 268 898 272
rect 870 258 874 262
rect 838 248 842 252
rect 830 168 834 172
rect 806 148 810 152
rect 878 158 882 162
rect 854 148 858 152
rect 870 148 874 152
rect 814 138 818 142
rect 846 138 850 142
rect 1126 658 1130 662
rect 1198 778 1202 782
rect 1158 748 1162 752
rect 1166 748 1170 752
rect 1222 818 1226 822
rect 1310 858 1314 862
rect 1326 838 1330 842
rect 1222 768 1226 772
rect 1190 738 1194 742
rect 1294 798 1298 802
rect 1246 768 1250 772
rect 1254 758 1258 762
rect 1230 748 1234 752
rect 1182 728 1186 732
rect 1166 708 1170 712
rect 1174 708 1178 712
rect 1158 658 1162 662
rect 1150 648 1154 652
rect 1174 658 1178 662
rect 1230 728 1234 732
rect 1246 688 1250 692
rect 1262 748 1266 752
rect 1262 728 1266 732
rect 1302 768 1306 772
rect 1318 768 1322 772
rect 1350 798 1354 802
rect 1366 748 1370 752
rect 1302 728 1306 732
rect 1382 778 1386 782
rect 1470 1088 1474 1092
rect 1462 1038 1466 1042
rect 1430 928 1434 932
rect 1446 928 1450 932
rect 1422 838 1426 842
rect 1454 838 1458 842
rect 1446 808 1450 812
rect 1446 778 1450 782
rect 1430 768 1434 772
rect 1414 758 1418 762
rect 1382 748 1386 752
rect 1398 748 1402 752
rect 1374 728 1378 732
rect 1342 718 1346 722
rect 1350 718 1354 722
rect 1374 718 1378 722
rect 1334 708 1338 712
rect 1366 708 1370 712
rect 1334 698 1338 702
rect 1358 688 1362 692
rect 1278 678 1282 682
rect 1334 678 1338 682
rect 1230 668 1234 672
rect 1246 668 1250 672
rect 1254 668 1258 672
rect 1302 668 1306 672
rect 1326 668 1330 672
rect 1206 658 1210 662
rect 1398 728 1402 732
rect 1422 748 1426 752
rect 1438 738 1442 742
rect 1382 678 1386 682
rect 1390 678 1394 682
rect 1398 678 1402 682
rect 1254 658 1258 662
rect 1286 658 1290 662
rect 1334 658 1338 662
rect 1358 658 1362 662
rect 1382 658 1386 662
rect 1406 658 1410 662
rect 1182 648 1186 652
rect 1302 648 1306 652
rect 1334 648 1338 652
rect 1110 638 1114 642
rect 1166 638 1170 642
rect 1206 638 1210 642
rect 1102 628 1106 632
rect 1198 618 1202 622
rect 1102 608 1106 612
rect 1126 598 1130 602
rect 1086 518 1090 522
rect 1030 408 1034 412
rect 1006 378 1010 382
rect 1054 378 1058 382
rect 1062 378 1066 382
rect 1022 358 1026 362
rect 1046 358 1050 362
rect 990 348 994 352
rect 1006 348 1010 352
rect 1078 468 1082 472
rect 1070 368 1074 372
rect 1038 348 1042 352
rect 1062 348 1066 352
rect 998 338 1002 342
rect 934 288 938 292
rect 1022 328 1026 332
rect 1054 328 1058 332
rect 976 303 980 307
rect 981 303 985 307
rect 986 303 990 307
rect 982 288 986 292
rect 966 278 970 282
rect 942 268 946 272
rect 942 178 946 182
rect 1086 438 1090 442
rect 1118 528 1122 532
rect 1134 578 1138 582
rect 1190 578 1194 582
rect 1190 568 1194 572
rect 1142 558 1146 562
rect 1134 548 1138 552
rect 1150 548 1154 552
rect 1142 518 1146 522
rect 1214 588 1218 592
rect 1294 638 1298 642
rect 1246 578 1250 582
rect 1254 578 1258 582
rect 1302 588 1306 592
rect 1230 568 1234 572
rect 1238 558 1242 562
rect 1302 558 1306 562
rect 1398 648 1402 652
rect 1398 578 1402 582
rect 1414 648 1418 652
rect 1454 768 1458 772
rect 1430 678 1434 682
rect 1422 598 1426 602
rect 1246 548 1250 552
rect 1278 548 1282 552
rect 1382 548 1386 552
rect 1406 548 1410 552
rect 1254 538 1258 542
rect 1270 538 1274 542
rect 1206 478 1210 482
rect 1182 458 1186 462
rect 1094 388 1098 392
rect 1110 368 1114 372
rect 1094 358 1098 362
rect 1102 358 1106 362
rect 1142 358 1146 362
rect 1126 348 1130 352
rect 1078 268 1082 272
rect 1030 258 1034 262
rect 1102 258 1106 262
rect 1054 238 1058 242
rect 1142 238 1146 242
rect 1006 158 1010 162
rect 1014 158 1018 162
rect 1014 148 1018 152
rect 894 138 898 142
rect 974 138 978 142
rect 1110 158 1114 162
rect 1062 148 1066 152
rect 1086 148 1090 152
rect 1102 148 1106 152
rect 1046 138 1050 142
rect 942 128 946 132
rect 958 128 962 132
rect 1022 128 1026 132
rect 862 118 866 122
rect 878 118 882 122
rect 798 88 802 92
rect 838 98 842 102
rect 806 78 810 82
rect 814 78 818 82
rect 976 103 980 107
rect 981 103 985 107
rect 986 103 990 107
rect 950 98 954 102
rect 1038 88 1042 92
rect 926 78 930 82
rect 934 78 938 82
rect 902 68 906 72
rect 750 58 754 62
rect 782 58 786 62
rect 1038 58 1042 62
rect 1070 108 1074 112
rect 1070 68 1074 72
rect 1214 468 1218 472
rect 1318 538 1322 542
rect 1318 528 1322 532
rect 1302 508 1306 512
rect 1270 488 1274 492
rect 1302 488 1306 492
rect 1294 468 1298 472
rect 1342 508 1346 512
rect 1358 508 1362 512
rect 1334 498 1338 502
rect 1246 458 1250 462
rect 1262 458 1266 462
rect 1278 458 1282 462
rect 1310 458 1314 462
rect 1214 388 1218 392
rect 1206 378 1210 382
rect 1158 358 1162 362
rect 1358 478 1362 482
rect 1374 518 1378 522
rect 1358 468 1362 472
rect 1406 488 1410 492
rect 1398 468 1402 472
rect 1486 998 1490 1002
rect 1486 858 1490 862
rect 1486 798 1490 802
rect 1478 738 1482 742
rect 1470 718 1474 722
rect 1446 588 1450 592
rect 1454 548 1458 552
rect 1438 538 1442 542
rect 1430 528 1434 532
rect 1454 528 1458 532
rect 1422 498 1426 502
rect 1486 698 1490 702
rect 1422 458 1426 462
rect 1406 448 1410 452
rect 1414 448 1418 452
rect 1398 438 1402 442
rect 1342 368 1346 372
rect 1222 358 1226 362
rect 1278 358 1282 362
rect 1350 358 1354 362
rect 1254 348 1258 352
rect 1286 348 1290 352
rect 1318 348 1322 352
rect 1334 348 1338 352
rect 1286 328 1290 332
rect 1238 318 1242 322
rect 1190 278 1194 282
rect 1430 388 1434 392
rect 1374 358 1378 362
rect 1486 358 1490 362
rect 1366 348 1370 352
rect 1366 338 1370 342
rect 1406 338 1410 342
rect 1334 288 1338 292
rect 1350 288 1354 292
rect 1358 288 1362 292
rect 1270 278 1274 282
rect 1302 278 1306 282
rect 1398 328 1402 332
rect 1414 328 1418 332
rect 1446 328 1450 332
rect 1438 318 1442 322
rect 1462 318 1466 322
rect 1390 288 1394 292
rect 1302 268 1306 272
rect 1158 258 1162 262
rect 1174 258 1178 262
rect 1270 258 1274 262
rect 1310 258 1314 262
rect 1326 258 1330 262
rect 1206 168 1210 172
rect 1214 158 1218 162
rect 1230 148 1234 152
rect 1102 128 1106 132
rect 1142 128 1146 132
rect 1286 148 1290 152
rect 1302 148 1306 152
rect 1454 278 1458 282
rect 1454 248 1458 252
rect 1438 148 1442 152
rect 1374 138 1378 142
rect 1318 118 1322 122
rect 1430 118 1434 122
rect 1486 258 1490 262
rect 1486 158 1490 162
rect 1446 78 1450 82
rect 1086 58 1090 62
rect 1134 58 1138 62
rect 1158 58 1162 62
rect 1182 58 1186 62
rect 1198 58 1202 62
rect 1214 58 1218 62
rect 1382 58 1386 62
rect 1406 58 1410 62
rect 1430 58 1434 62
rect 1462 58 1466 62
rect 742 38 746 42
rect 966 38 970 42
rect 998 38 1002 42
rect 1062 38 1066 42
rect 886 8 890 12
rect 918 8 922 12
rect 1022 8 1026 12
rect 1038 8 1042 12
<< metal3 >>
rect 874 1208 886 1211
rect 898 1208 910 1211
rect 922 1208 934 1211
rect 1042 1208 1054 1211
rect 1066 1208 1078 1211
rect 1242 1208 1254 1211
rect 166 1202 169 1208
rect 486 1203 488 1207
rect 614 1202 617 1208
rect 998 1202 1001 1208
rect 1106 1198 1118 1201
rect 1114 1188 1134 1191
rect 202 1168 214 1171
rect 218 1168 318 1171
rect 410 1158 422 1161
rect 658 1158 662 1161
rect 1490 1158 1513 1161
rect 70 1151 73 1158
rect 142 1151 145 1158
rect 70 1148 145 1151
rect 178 1148 390 1151
rect 442 1148 526 1151
rect 638 1151 641 1158
rect 734 1151 737 1158
rect 638 1148 737 1151
rect 858 1148 870 1151
rect 874 1148 894 1151
rect 1178 1148 1297 1151
rect 1418 1148 1438 1151
rect 1442 1148 1446 1151
rect 414 1141 417 1148
rect 1294 1142 1297 1148
rect 386 1138 417 1141
rect 678 1138 790 1141
rect 1082 1138 1094 1141
rect 1154 1138 1238 1141
rect 1298 1138 1398 1141
rect 10 1128 126 1131
rect 130 1128 174 1131
rect 370 1128 446 1131
rect 454 1131 457 1138
rect 678 1132 681 1138
rect 454 1128 558 1131
rect 674 1128 678 1131
rect 190 1121 193 1128
rect 190 1118 406 1121
rect 410 1118 518 1121
rect 554 1118 582 1121
rect 586 1118 598 1121
rect 978 1118 1014 1121
rect 166 1112 169 1118
rect 290 1108 334 1111
rect 378 1108 430 1111
rect 546 1108 630 1111
rect 754 1108 782 1111
rect 786 1108 878 1111
rect 1050 1108 1062 1111
rect 1090 1108 1142 1111
rect 990 1103 992 1107
rect 1026 1098 1070 1101
rect 1098 1098 1134 1101
rect 682 1088 686 1091
rect 690 1088 742 1091
rect 890 1088 926 1091
rect 930 1088 950 1091
rect 954 1088 1078 1091
rect 1298 1088 1342 1091
rect 1362 1088 1406 1091
rect 1410 1088 1470 1091
rect 62 1078 129 1081
rect 62 1072 65 1078
rect 126 1072 129 1078
rect 402 1078 462 1081
rect 530 1078 670 1081
rect 1086 1081 1089 1088
rect 1086 1078 1166 1081
rect 1210 1078 1246 1081
rect 1382 1078 1390 1081
rect 286 1071 289 1078
rect 1382 1072 1385 1078
rect 202 1068 374 1071
rect 414 1068 470 1071
rect 474 1068 510 1071
rect 562 1068 582 1071
rect 586 1068 614 1071
rect 930 1068 993 1071
rect 1058 1068 1126 1071
rect 1170 1068 1222 1071
rect 1290 1068 1310 1071
rect 414 1062 417 1068
rect 990 1062 993 1068
rect -26 1058 6 1061
rect 90 1058 142 1061
rect 254 1058 289 1061
rect 434 1058 454 1061
rect 594 1058 622 1061
rect 626 1058 654 1061
rect 726 1058 798 1061
rect 1138 1058 1166 1061
rect 1170 1058 1294 1061
rect 1298 1058 1350 1061
rect 1378 1058 1414 1061
rect 254 1052 257 1058
rect 286 1052 289 1058
rect 442 1048 566 1051
rect 570 1048 590 1051
rect 642 1048 646 1051
rect 670 1051 673 1058
rect 726 1052 729 1058
rect 670 1048 678 1051
rect 970 1048 1094 1051
rect 1098 1048 1174 1051
rect 1210 1048 1214 1051
rect 1218 1048 1270 1051
rect 1274 1048 1318 1051
rect 1322 1048 1358 1051
rect 614 1042 617 1048
rect 338 1038 446 1041
rect 1210 1038 1289 1041
rect 1306 1038 1462 1041
rect 1286 1032 1289 1038
rect 998 1012 1001 1018
rect 486 1003 488 1007
rect 690 998 814 1001
rect 818 998 846 1001
rect 1490 998 1513 1001
rect 6 981 9 988
rect -26 978 9 981
rect 1338 978 1398 981
rect 1422 981 1425 988
rect 1422 978 1513 981
rect 26 968 142 971
rect 146 968 190 971
rect 194 968 246 971
rect 402 968 430 971
rect 594 968 649 971
rect 906 968 1110 971
rect 1162 968 1190 971
rect 1254 971 1257 978
rect 1242 968 1257 971
rect 1378 968 1406 971
rect 646 962 649 968
rect -26 958 30 961
rect 322 958 438 961
rect 578 958 630 961
rect 1178 958 1190 961
rect 1194 958 1366 961
rect 1442 958 1513 961
rect 214 951 217 958
rect 262 951 265 958
rect 214 948 265 951
rect 322 948 326 951
rect 362 948 454 951
rect 458 948 510 951
rect 554 948 622 951
rect 634 948 678 951
rect 750 951 753 958
rect 714 948 753 951
rect 910 951 913 958
rect 910 948 942 951
rect 946 948 1150 951
rect 1170 948 1214 951
rect 1266 948 1398 951
rect 134 941 137 948
rect 134 938 182 941
rect 294 941 297 948
rect 294 938 326 941
rect 358 938 430 941
rect 682 938 822 941
rect 858 938 862 941
rect 866 938 894 941
rect 898 938 918 941
rect 1126 938 1134 941
rect 1138 938 1238 941
rect 1274 938 1382 941
rect 1430 941 1433 948
rect 1390 938 1433 941
rect 358 932 361 938
rect 526 931 529 938
rect 410 928 529 931
rect 558 931 561 938
rect 1390 932 1393 938
rect 558 928 574 931
rect 626 928 702 931
rect 978 928 1254 931
rect 1434 928 1446 931
rect 122 918 142 921
rect 274 918 302 921
rect 418 918 534 921
rect 538 918 582 921
rect 970 918 1174 921
rect 1238 918 1246 921
rect 1250 918 1302 921
rect 250 908 334 911
rect 1034 908 1054 911
rect 1154 908 1166 911
rect 990 903 992 907
rect 154 898 158 901
rect 162 898 718 901
rect 722 898 726 901
rect 1130 898 1142 901
rect 1146 898 1214 901
rect 50 888 286 891
rect 290 888 462 891
rect 466 888 534 891
rect 538 888 566 891
rect 574 888 622 891
rect 754 888 838 891
rect 874 888 878 891
rect 1090 888 1150 891
rect 574 881 577 888
rect 514 878 577 881
rect 602 878 646 881
rect 650 878 774 881
rect 786 878 862 881
rect 938 878 950 881
rect 126 871 129 878
rect 66 868 129 871
rect 178 868 185 871
rect 350 871 353 878
rect 234 868 353 871
rect 358 868 470 871
rect 650 868 654 871
rect 698 868 718 871
rect 862 871 865 878
rect 862 868 950 871
rect 1074 868 1094 871
rect 1194 868 1198 871
rect 182 862 185 868
rect -26 858 6 861
rect 186 858 246 861
rect 358 861 361 868
rect 338 858 361 861
rect 434 858 446 861
rect 490 858 542 861
rect 574 861 577 868
rect 574 858 582 861
rect 610 858 630 861
rect 746 858 878 861
rect 946 858 1014 861
rect 1078 858 1086 861
rect 1090 858 1102 861
rect 1106 858 1190 861
rect 1194 858 1310 861
rect 1490 858 1513 861
rect 218 848 278 851
rect 458 848 494 851
rect 570 848 582 851
rect 594 848 654 851
rect 826 848 958 851
rect 962 848 982 851
rect 1106 848 1166 851
rect 98 838 310 841
rect 346 838 438 841
rect 538 838 686 841
rect 938 838 1070 841
rect 1090 838 1142 841
rect 1202 838 1206 841
rect 1210 838 1326 841
rect 1330 838 1422 841
rect 1426 838 1454 841
rect 138 828 190 831
rect 442 828 478 831
rect 482 828 518 831
rect 874 828 990 831
rect 1002 828 1182 831
rect 202 818 222 821
rect 226 818 942 821
rect 1066 818 1222 821
rect 714 808 718 811
rect 730 808 878 811
rect 882 808 1438 811
rect 1442 808 1446 811
rect 486 803 488 807
rect 1098 798 1126 801
rect 1298 798 1350 801
rect 1490 798 1513 801
rect 626 788 702 791
rect 706 788 830 791
rect 994 788 1102 791
rect 362 778 510 781
rect 578 778 678 781
rect 778 778 790 781
rect 794 778 830 781
rect 834 778 1038 781
rect 1090 778 1126 781
rect 1154 778 1198 781
rect 1450 778 1513 781
rect 130 768 246 771
rect 410 768 598 771
rect 898 768 974 771
rect 986 768 990 771
rect 994 768 1070 771
rect 1142 771 1145 778
rect 1142 768 1222 771
rect 1250 768 1302 771
rect 1382 771 1385 778
rect 1322 768 1385 771
rect 1434 768 1454 771
rect -26 758 6 761
rect 162 758 166 761
rect 170 758 254 761
rect 390 761 393 768
rect 390 758 462 761
rect 698 758 798 761
rect 814 761 817 768
rect 814 758 854 761
rect 858 758 886 761
rect 914 758 1038 761
rect 1122 758 1158 761
rect 1170 758 1254 761
rect 1366 758 1374 761
rect 1418 758 1513 761
rect 74 748 134 751
rect 294 748 302 751
rect 310 751 313 758
rect 1366 752 1369 758
rect 310 748 422 751
rect 522 748 566 751
rect 570 748 662 751
rect 850 748 886 751
rect 914 748 1134 751
rect 1138 748 1158 751
rect 1162 748 1166 751
rect 1234 748 1262 751
rect 1386 748 1398 751
rect 1402 748 1422 751
rect 66 738 118 741
rect 122 738 182 741
rect 242 738 278 741
rect 378 738 398 741
rect 434 738 462 741
rect 506 738 550 741
rect 898 738 918 741
rect 1010 738 1014 741
rect 1042 738 1190 741
rect 1194 738 1438 741
rect 1482 738 1513 741
rect 42 728 54 731
rect 98 728 158 731
rect 210 728 230 731
rect 250 728 254 731
rect 278 731 281 738
rect 278 728 286 731
rect 290 728 294 731
rect 298 728 310 731
rect 370 728 398 731
rect 458 728 542 731
rect 794 728 814 731
rect 970 728 1086 731
rect 1090 728 1142 731
rect 1162 728 1182 731
rect 1234 728 1262 731
rect 1306 728 1374 731
rect 1378 728 1398 731
rect 106 718 126 721
rect 258 718 318 721
rect 322 718 326 721
rect 330 718 382 721
rect 490 718 518 721
rect 714 718 726 721
rect 818 718 942 721
rect 946 718 966 721
rect 978 718 1134 721
rect 1274 718 1342 721
rect 1354 718 1374 721
rect 1474 718 1513 721
rect 730 708 910 711
rect 1058 708 1166 711
rect 1178 708 1278 711
rect 1338 708 1366 711
rect 990 703 992 707
rect 178 698 206 701
rect 546 698 590 701
rect 770 698 806 701
rect 810 698 830 701
rect 834 698 846 701
rect 866 698 953 701
rect 1098 698 1126 701
rect 1130 698 1334 701
rect 1490 698 1513 701
rect 74 688 254 691
rect 258 688 270 691
rect 554 688 606 691
rect 874 688 902 691
rect 914 688 942 691
rect 950 691 953 698
rect 950 688 1006 691
rect 1362 688 1393 691
rect 194 678 222 681
rect 434 678 542 681
rect 546 678 702 681
rect 842 678 862 681
rect 866 678 1054 681
rect 1246 681 1249 688
rect 1390 682 1393 688
rect 1246 678 1278 681
rect 1338 678 1382 681
rect 1434 678 1513 681
rect 126 671 129 678
rect 42 668 129 671
rect 146 668 278 671
rect 282 668 326 671
rect 338 668 374 671
rect 402 668 414 671
rect 418 668 430 671
rect 626 668 646 671
rect 702 668 705 678
rect 794 668 822 671
rect 826 668 846 671
rect 850 668 894 671
rect 906 668 926 671
rect 1122 668 1230 671
rect 1250 668 1254 671
rect 1258 668 1302 671
rect 1398 671 1401 678
rect 1330 668 1401 671
rect -26 658 6 661
rect 94 658 161 661
rect 210 658 254 661
rect 258 658 358 661
rect 410 658 550 661
rect 706 658 710 661
rect 818 658 854 661
rect 858 658 902 661
rect 958 661 961 668
rect 958 658 1054 661
rect 1130 658 1158 661
rect 1210 658 1254 661
rect 1258 658 1270 661
rect 1278 658 1286 661
rect 1338 658 1358 661
rect 1386 658 1406 661
rect 1490 658 1513 661
rect 94 652 97 658
rect 158 652 161 658
rect 374 648 382 651
rect 386 648 430 651
rect 490 648 574 651
rect 578 648 598 651
rect 602 648 633 651
rect 778 648 870 651
rect 970 648 1078 651
rect 1094 651 1097 658
rect 1094 648 1102 651
rect 1174 651 1177 658
rect 1154 648 1177 651
rect 1186 648 1193 651
rect 1306 648 1334 651
rect 1338 648 1345 651
rect 1402 648 1414 651
rect 274 638 334 641
rect 350 641 353 648
rect 630 642 633 648
rect 350 638 470 641
rect 474 638 534 641
rect 538 638 558 641
rect 1066 638 1110 641
rect 1170 638 1206 641
rect 1298 638 1486 641
rect 946 628 966 631
rect 1082 628 1102 631
rect 1106 628 1201 631
rect 1198 622 1201 628
rect 394 618 726 621
rect 786 618 846 621
rect 722 608 782 611
rect 1106 608 1214 611
rect 486 603 488 607
rect 970 598 1038 601
rect 1042 598 1126 601
rect 1426 598 1513 601
rect 66 588 86 591
rect 90 588 190 591
rect 314 588 398 591
rect 1034 588 1193 591
rect 1218 588 1302 591
rect 6 581 9 588
rect -26 578 9 581
rect 298 578 342 581
rect 346 578 542 581
rect 878 581 881 588
rect 1190 582 1193 588
rect 878 578 918 581
rect 1242 578 1246 581
rect 1446 581 1449 588
rect 1446 578 1513 581
rect 850 568 942 571
rect 1134 571 1137 578
rect 1134 568 1190 571
rect 1254 571 1257 578
rect 1234 568 1257 571
rect 1398 571 1401 578
rect 1398 568 1513 571
rect -26 558 30 561
rect 242 558 414 561
rect 582 561 585 568
rect 418 558 585 561
rect 906 558 910 561
rect 930 558 1014 561
rect 1138 558 1142 561
rect 1242 558 1302 561
rect 1510 558 1513 568
rect 58 548 94 551
rect 98 548 126 551
rect 158 551 161 558
rect 158 548 214 551
rect 354 548 366 551
rect 442 548 470 551
rect 554 548 646 551
rect 650 548 694 551
rect 714 548 822 551
rect 866 548 902 551
rect 1138 548 1150 551
rect 1154 548 1246 551
rect 1282 548 1382 551
rect 1386 548 1406 551
rect 1410 548 1446 551
rect 1450 548 1454 551
rect 178 538 257 541
rect 422 541 425 548
rect 410 538 425 541
rect 434 538 542 541
rect 610 538 638 541
rect 690 538 702 541
rect 762 538 1254 541
rect 1258 538 1270 541
rect 1322 538 1438 541
rect 254 532 257 538
rect 10 528 22 531
rect 26 528 46 531
rect 402 528 494 531
rect 658 528 742 531
rect 770 528 910 531
rect 930 528 934 531
rect 1010 528 1118 531
rect 1122 528 1246 531
rect 1250 528 1318 531
rect 1434 528 1454 531
rect 234 518 270 521
rect 306 518 630 521
rect 634 518 718 521
rect 722 518 726 521
rect 730 518 774 521
rect 802 518 814 521
rect 826 518 870 521
rect 898 518 902 521
rect 910 518 1086 521
rect 1090 518 1142 521
rect 1510 521 1513 531
rect 1378 518 1513 521
rect 370 508 422 511
rect 910 511 913 518
rect 834 508 913 511
rect 1026 508 1302 511
rect 1306 508 1342 511
rect 1346 508 1358 511
rect 990 503 992 507
rect 186 498 254 501
rect 258 498 310 501
rect 314 498 646 501
rect 650 498 694 501
rect 810 498 830 501
rect 842 498 894 501
rect 1338 498 1422 501
rect 66 488 102 491
rect 794 488 822 491
rect 842 488 910 491
rect 938 488 942 491
rect 1274 488 1302 491
rect 1306 488 1406 491
rect 90 478 174 481
rect 250 478 286 481
rect 290 478 614 481
rect 618 478 630 481
rect 634 478 654 481
rect 658 478 670 481
rect 734 481 737 488
rect 714 478 737 481
rect 762 478 1014 481
rect 1210 478 1358 481
rect 74 468 102 471
rect 122 468 150 471
rect 154 468 158 471
rect 210 468 342 471
rect 650 468 750 471
rect 882 468 886 471
rect 914 468 966 471
rect 1082 468 1185 471
rect 1218 468 1294 471
rect 1362 468 1398 471
rect 198 461 201 468
rect -26 458 206 461
rect 258 458 334 461
rect 430 458 446 461
rect 758 461 761 468
rect 738 458 761 461
rect 902 461 905 468
rect 1182 462 1185 468
rect 866 458 905 461
rect 914 458 998 461
rect 1250 458 1262 461
rect 1282 458 1310 461
rect 1426 458 1513 461
rect 430 452 433 458
rect 130 448 166 451
rect 170 448 206 451
rect 454 448 566 451
rect 570 448 638 451
rect 686 451 689 458
rect 686 448 774 451
rect 802 448 838 451
rect 842 448 894 451
rect 930 448 934 451
rect 954 448 958 451
rect 1410 448 1414 451
rect 194 438 262 441
rect 278 441 281 448
rect 266 438 281 441
rect 298 438 342 441
rect 454 441 457 448
rect 346 438 457 441
rect 578 438 598 441
rect 746 438 814 441
rect 886 438 918 441
rect 926 438 942 441
rect 958 438 1086 441
rect 1386 438 1398 441
rect 886 432 889 438
rect 926 432 929 438
rect 958 432 961 438
rect 538 418 942 421
rect 1030 412 1033 421
rect 486 403 488 407
rect 362 388 526 391
rect 554 388 766 391
rect 778 388 910 391
rect 1098 388 1214 391
rect 138 378 238 381
rect 346 378 582 381
rect 634 378 670 381
rect 674 378 798 381
rect 1010 378 1054 381
rect 1066 378 1206 381
rect 1430 381 1433 388
rect 1430 378 1513 381
rect 234 368 257 371
rect 254 362 257 368
rect 618 368 630 371
rect 730 368 750 371
rect 778 368 790 371
rect 802 368 830 371
rect 834 368 1070 371
rect 1114 368 1342 371
rect -26 358 6 361
rect 330 358 374 361
rect 406 361 409 368
rect 378 358 409 361
rect 522 358 846 361
rect 898 358 1022 361
rect 1038 358 1046 361
rect 1050 358 1094 361
rect 1106 358 1142 361
rect 1162 358 1222 361
rect 1226 358 1278 361
rect 1282 358 1350 361
rect 1354 358 1374 361
rect 1490 358 1513 361
rect 94 351 97 358
rect 94 348 142 351
rect 202 348 222 351
rect 278 351 281 358
rect 274 348 281 351
rect 290 348 342 351
rect 402 348 462 351
rect 482 348 534 351
rect 586 348 606 351
rect 698 348 742 351
rect 746 348 766 351
rect 786 348 894 351
rect 994 348 1006 351
rect 1042 348 1062 351
rect 1290 348 1318 351
rect 1338 348 1366 351
rect 178 338 214 341
rect 218 338 302 341
rect 442 338 558 341
rect 642 338 758 341
rect 762 338 878 341
rect 1002 338 1070 341
rect 1126 341 1129 348
rect 1254 341 1257 348
rect 1406 342 1409 348
rect 1074 338 1366 341
rect 62 331 65 338
rect 126 331 129 338
rect 62 328 129 331
rect 290 328 326 331
rect 366 331 369 338
rect 366 328 438 331
rect 458 328 518 331
rect 522 328 574 331
rect 602 328 662 331
rect 682 328 686 331
rect 690 328 710 331
rect 866 328 878 331
rect 1026 328 1054 331
rect 1238 328 1286 331
rect 1402 328 1414 331
rect 1418 328 1446 331
rect 1238 322 1241 328
rect 178 318 422 321
rect 434 318 598 321
rect 610 318 678 321
rect 1442 318 1462 321
rect 314 308 374 311
rect 466 308 534 311
rect 538 308 694 311
rect 990 303 992 307
rect 10 298 246 301
rect 322 298 462 301
rect 522 298 726 301
rect 210 288 270 291
rect 394 288 398 291
rect 642 288 814 291
rect 938 288 982 291
rect 1338 288 1350 291
rect 1362 288 1390 291
rect 202 278 414 281
rect 442 278 510 281
rect 514 278 518 281
rect 546 278 598 281
rect 658 278 758 281
rect 770 278 798 281
rect 802 278 966 281
rect 1274 278 1302 281
rect 1306 278 1454 281
rect 202 268 209 271
rect 70 261 73 268
rect 206 262 209 268
rect 362 268 382 271
rect 426 268 446 271
rect 458 268 542 271
rect 586 268 590 271
rect 722 268 854 271
rect 858 268 894 271
rect 946 268 1078 271
rect 1190 271 1193 278
rect 1082 268 1193 271
rect 1274 268 1302 271
rect 70 258 78 261
rect 106 258 174 261
rect 310 261 313 268
rect 310 258 446 261
rect 506 258 521 261
rect 530 258 550 261
rect 574 261 577 268
rect 570 258 577 261
rect 642 258 654 261
rect 762 258 814 261
rect 874 258 902 261
rect 906 258 1030 261
rect 1106 258 1158 261
rect 1178 258 1270 261
rect 1274 258 1310 261
rect 1314 258 1326 261
rect 1490 258 1513 261
rect 518 252 521 258
rect 122 248 126 251
rect 194 248 398 251
rect 402 248 414 251
rect 586 248 598 251
rect 614 251 617 258
rect 614 248 686 251
rect 822 251 825 258
rect 794 248 838 251
rect 1370 248 1454 251
rect 250 238 326 241
rect 482 238 494 241
rect 550 238 558 241
rect 578 238 614 241
rect 634 238 646 241
rect 1058 238 1142 241
rect 654 232 657 238
rect 314 228 478 231
rect 490 228 550 231
rect 274 218 486 221
rect 646 212 649 221
rect 486 203 488 207
rect 494 198 654 201
rect 658 198 774 201
rect 114 188 166 191
rect 170 188 278 191
rect 494 191 497 198
rect 330 188 497 191
rect 522 188 590 191
rect 642 188 654 191
rect 210 178 286 181
rect 522 178 526 181
rect 694 181 697 188
rect 554 178 697 181
rect 754 178 942 181
rect 114 168 134 171
rect 138 168 254 171
rect 258 168 302 171
rect 426 168 558 171
rect 594 168 606 171
rect 634 168 830 171
rect 1210 168 1438 171
rect 266 158 310 161
rect 394 158 398 161
rect 402 158 430 161
rect 434 158 454 161
rect 458 158 478 161
rect 574 161 577 168
rect 546 158 662 161
rect 882 158 1006 161
rect 1018 158 1022 161
rect 1106 158 1110 161
rect 1490 158 1513 161
rect 134 151 137 158
rect 90 148 137 151
rect 166 151 169 158
rect 198 151 201 158
rect 286 152 289 158
rect 166 148 201 151
rect 226 148 249 151
rect 354 148 374 151
rect 402 148 638 151
rect 650 148 654 151
rect 722 148 729 151
rect 810 148 854 151
rect 874 148 881 151
rect 1018 148 1062 151
rect 1066 148 1086 151
rect 1090 148 1102 151
rect 1214 151 1217 158
rect 1438 152 1441 158
rect 1106 148 1217 151
rect 1234 148 1286 151
rect 1306 148 1377 151
rect 210 138 238 141
rect 246 141 249 148
rect 1374 142 1377 148
rect 246 138 318 141
rect 370 138 414 141
rect 418 138 470 141
rect 474 138 614 141
rect 618 138 622 141
rect 626 138 678 141
rect 690 138 694 141
rect 714 138 734 141
rect 818 138 846 141
rect 898 138 974 141
rect 1042 138 1046 141
rect 66 128 214 131
rect 370 128 454 131
rect 530 128 598 131
rect 706 128 782 131
rect 946 128 958 131
rect 1106 128 1142 131
rect 518 122 521 128
rect 18 118 22 121
rect 170 118 206 121
rect 274 118 510 121
rect 554 118 558 121
rect 754 118 862 121
rect 866 118 873 121
rect 1022 121 1025 128
rect 882 118 1025 121
rect 1322 118 1430 121
rect 1070 112 1073 118
rect 98 108 182 111
rect 242 108 366 111
rect 370 108 398 111
rect 410 108 430 111
rect 498 108 510 111
rect 990 103 992 107
rect 186 98 238 101
rect 354 98 438 101
rect 482 98 566 101
rect 570 98 718 101
rect 842 98 950 101
rect 74 88 118 91
rect 162 88 222 91
rect 298 88 382 91
rect 418 88 470 91
rect 714 88 798 91
rect 934 88 1038 91
rect -26 78 30 81
rect 90 78 102 81
rect 106 78 158 81
rect 210 78 358 81
rect 362 78 422 81
rect 534 78 537 88
rect 934 82 937 88
rect 554 78 806 81
rect 818 78 926 81
rect 42 68 89 71
rect 122 68 126 71
rect 130 68 286 71
rect 290 68 294 71
rect 442 68 486 71
rect 514 68 582 71
rect 782 68 902 71
rect 1446 68 1449 78
rect -26 58 6 61
rect 58 58 78 61
rect 86 61 89 68
rect 86 58 182 61
rect 186 58 230 61
rect 298 58 326 61
rect 330 58 422 61
rect 462 58 534 61
rect 626 58 670 61
rect 694 61 697 68
rect 782 62 785 68
rect 694 58 750 61
rect 902 61 905 68
rect 902 58 1038 61
rect 1070 61 1073 68
rect 1070 58 1086 61
rect 1138 58 1158 61
rect 1162 58 1182 61
rect 1186 58 1198 61
rect 1202 58 1214 61
rect 1386 58 1406 61
rect 1410 58 1430 61
rect 1434 58 1462 61
rect 462 52 465 58
rect 162 48 190 51
rect 258 48 438 51
rect 510 48 518 51
rect 522 48 582 51
rect 642 48 662 51
rect 314 38 622 41
rect 698 38 742 41
rect 970 38 998 41
rect 1002 38 1062 41
rect 590 12 593 18
rect 886 12 889 18
rect 1038 12 1041 18
rect 626 8 630 11
rect 922 8 926 11
rect 1018 8 1022 11
rect 486 3 488 7
<< m4contact >>
rect 473 1203 476 1207
rect 476 1203 477 1207
rect 479 1203 481 1207
rect 481 1203 482 1207
rect 482 1203 483 1207
rect 166 1198 170 1202
rect 614 1198 618 1202
rect 998 1198 1002 1202
rect 670 1128 674 1132
rect 166 1118 170 1122
rect 977 1103 980 1107
rect 980 1103 981 1107
rect 983 1103 985 1107
rect 985 1103 986 1107
rect 986 1103 987 1107
rect 886 1088 890 1092
rect 1406 1088 1410 1092
rect 1390 1078 1394 1082
rect 1350 1058 1354 1062
rect 614 1048 618 1052
rect 678 1048 682 1052
rect 1206 1048 1210 1052
rect 998 1018 1002 1022
rect 473 1003 476 1007
rect 476 1003 477 1007
rect 479 1003 481 1007
rect 481 1003 482 1007
rect 482 1003 483 1007
rect 977 903 980 907
rect 980 903 981 907
rect 983 903 985 907
rect 985 903 986 907
rect 986 903 987 907
rect 150 898 154 902
rect 726 898 730 902
rect 1126 898 1130 902
rect 870 888 874 892
rect 934 878 938 882
rect 174 868 178 872
rect 878 858 882 862
rect 1190 858 1194 862
rect 198 818 202 822
rect 710 808 714 812
rect 726 808 730 812
rect 1438 808 1442 812
rect 473 803 476 807
rect 476 803 477 807
rect 479 803 481 807
rect 481 803 482 807
rect 482 803 483 807
rect 1126 798 1130 802
rect 702 788 706 792
rect 1126 778 1130 782
rect 1150 778 1154 782
rect 974 768 978 772
rect 1158 758 1162 762
rect 1374 758 1378 762
rect 302 748 306 752
rect 182 738 186 742
rect 1006 738 1010 742
rect 1158 728 1162 732
rect 966 718 970 722
rect 974 718 978 722
rect 1270 718 1274 722
rect 1350 718 1354 722
rect 1278 708 1282 712
rect 977 703 980 707
rect 980 703 981 707
rect 983 703 985 707
rect 985 703 986 707
rect 986 703 987 707
rect 1094 698 1098 702
rect 902 688 906 692
rect 702 678 706 682
rect 430 668 434 672
rect 894 668 898 672
rect 902 668 906 672
rect 710 658 714 662
rect 1270 658 1274 662
rect 1286 658 1290 662
rect 1486 658 1490 662
rect 966 648 970 652
rect 1102 648 1106 652
rect 1182 648 1186 652
rect 1486 638 1490 642
rect 726 618 730 622
rect 718 608 722 612
rect 1214 608 1218 612
rect 473 603 476 607
rect 476 603 477 607
rect 479 603 481 607
rect 481 603 482 607
rect 482 603 483 607
rect 294 578 298 582
rect 1238 578 1242 582
rect 910 558 914 562
rect 1014 558 1018 562
rect 1134 558 1138 562
rect 1446 548 1450 552
rect 430 538 434 542
rect 926 528 930 532
rect 1246 528 1250 532
rect 894 518 898 522
rect 977 503 980 507
rect 980 503 981 507
rect 983 503 985 507
rect 985 503 986 507
rect 986 503 987 507
rect 894 498 898 502
rect 910 488 914 492
rect 942 488 946 492
rect 150 468 154 472
rect 750 468 754 472
rect 886 468 890 472
rect 910 468 914 472
rect 206 458 210 462
rect 926 448 930 452
rect 950 448 954 452
rect 294 438 298 442
rect 918 438 922 442
rect 1382 438 1386 442
rect 1030 408 1034 412
rect 473 403 476 407
rect 476 403 477 407
rect 479 403 481 407
rect 481 403 482 407
rect 482 403 483 407
rect 630 368 634 372
rect 894 358 898 362
rect 270 348 274 352
rect 478 348 482 352
rect 1006 348 1010 352
rect 1406 348 1410 352
rect 1070 338 1074 342
rect 534 308 538 312
rect 977 303 980 307
rect 980 303 981 307
rect 983 303 985 307
rect 985 303 986 307
rect 986 303 987 307
rect 398 288 402 292
rect 638 288 642 292
rect 518 278 522 282
rect 198 268 202 272
rect 454 268 458 272
rect 582 268 586 272
rect 1270 268 1274 272
rect 78 258 82 262
rect 550 258 554 262
rect 654 258 658 262
rect 902 258 906 262
rect 1030 258 1034 262
rect 126 248 130 252
rect 414 248 418 252
rect 1366 248 1370 252
rect 558 238 562 242
rect 646 238 650 242
rect 654 228 658 232
rect 646 208 650 212
rect 473 203 476 207
rect 476 203 477 207
rect 479 203 481 207
rect 481 203 482 207
rect 482 203 483 207
rect 654 188 658 192
rect 518 178 522 182
rect 750 178 754 182
rect 1438 168 1442 172
rect 390 158 394 162
rect 1022 158 1026 162
rect 1102 158 1106 162
rect 1438 158 1442 162
rect 398 148 402 152
rect 646 148 650 152
rect 718 148 722 152
rect 870 148 874 152
rect 694 138 698 142
rect 1038 138 1042 142
rect 518 128 522 132
rect 206 118 210 122
rect 510 118 514 122
rect 550 118 554 122
rect 1070 118 1074 122
rect 398 108 402 112
rect 977 103 980 107
rect 980 103 981 107
rect 983 103 985 107
rect 985 103 986 107
rect 986 103 987 107
rect 414 88 418 92
rect 534 88 538 92
rect 1446 78 1450 82
rect 118 68 122 72
rect 294 68 298 72
rect 510 68 514 72
rect 590 18 594 22
rect 886 18 890 22
rect 1038 18 1042 22
rect 622 8 626 12
rect 926 8 930 12
rect 1014 8 1018 12
rect 473 3 476 7
rect 476 3 477 7
rect 479 3 481 7
rect 481 3 482 7
rect 482 3 483 7
<< metal4 >>
rect 486 1203 488 1207
rect 166 1122 169 1198
rect 614 1052 617 1198
rect 670 1051 673 1128
rect 990 1103 992 1107
rect 670 1048 678 1051
rect 486 1003 488 1007
rect 718 898 726 901
rect 150 472 153 898
rect 178 868 185 871
rect 182 742 185 868
rect 198 461 201 818
rect 486 803 488 807
rect 294 748 302 751
rect 294 582 297 748
rect 702 682 705 788
rect 430 542 433 668
rect 710 662 713 808
rect 718 612 721 898
rect 874 888 881 891
rect 878 862 881 888
rect 726 622 729 808
rect 886 671 889 1088
rect 998 1022 1001 1198
rect 1382 1078 1390 1081
rect 1210 1048 1217 1051
rect 990 903 992 907
rect 902 672 905 688
rect 886 668 894 671
rect 486 603 488 607
rect 902 558 910 561
rect 894 522 897 528
rect 198 458 206 461
rect 274 348 286 351
rect 202 268 209 271
rect 70 258 78 261
rect 118 248 126 251
rect 118 72 121 248
rect 206 122 209 268
rect 294 72 297 438
rect 486 403 488 407
rect 474 348 478 351
rect 390 288 398 291
rect 390 162 393 288
rect 454 262 457 268
rect 398 112 401 148
rect 414 92 417 248
rect 486 203 488 207
rect 518 182 521 278
rect 518 132 521 148
rect 510 72 513 118
rect 534 92 537 308
rect 586 268 593 271
rect 554 258 558 261
rect 550 238 558 241
rect 550 122 553 238
rect 590 22 593 268
rect 630 11 633 368
rect 638 241 641 288
rect 646 258 654 261
rect 646 252 649 258
rect 638 238 646 241
rect 646 152 649 208
rect 654 192 657 228
rect 750 182 753 468
rect 722 148 729 151
rect 874 148 881 151
rect 878 142 881 148
rect 698 138 702 141
rect 886 22 889 468
rect 894 362 897 498
rect 902 262 905 558
rect 922 528 926 531
rect 934 491 937 878
rect 1126 802 1129 898
rect 1130 778 1134 781
rect 1146 778 1150 781
rect 974 722 977 768
rect 966 652 969 718
rect 990 703 992 707
rect 990 503 992 507
rect 934 488 942 491
rect 910 472 913 488
rect 954 448 961 451
rect 918 442 921 448
rect 626 8 633 11
rect 926 12 929 448
rect 1006 352 1009 738
rect 1158 732 1161 758
rect 1094 651 1097 698
rect 1094 648 1102 651
rect 1190 651 1193 858
rect 1186 648 1193 651
rect 1018 558 1022 561
rect 990 303 992 307
rect 1030 262 1033 408
rect 990 103 992 107
rect 1022 11 1025 158
rect 1038 22 1041 138
rect 1070 122 1073 338
rect 1102 162 1105 648
rect 1214 612 1217 1048
rect 1350 722 1353 1058
rect 1366 758 1374 761
rect 1270 662 1273 718
rect 1278 661 1281 708
rect 1278 658 1286 661
rect 1242 578 1249 581
rect 1138 558 1145 561
rect 1246 532 1249 578
rect 1270 272 1273 658
rect 1366 252 1369 758
rect 1382 442 1385 1078
rect 1406 352 1409 1088
rect 1438 172 1441 808
rect 1486 642 1489 658
rect 1438 162 1441 168
rect 1446 82 1449 548
rect 1018 8 1025 11
rect 486 3 488 7
<< m5contact >>
rect 472 1203 473 1207
rect 473 1203 476 1207
rect 477 1203 479 1207
rect 479 1203 481 1207
rect 482 1203 483 1207
rect 483 1203 486 1207
rect 976 1103 977 1107
rect 977 1103 980 1107
rect 981 1103 983 1107
rect 983 1103 985 1107
rect 986 1103 987 1107
rect 987 1103 990 1107
rect 472 1003 473 1007
rect 473 1003 476 1007
rect 477 1003 479 1007
rect 479 1003 481 1007
rect 482 1003 483 1007
rect 483 1003 486 1007
rect 472 803 473 807
rect 473 803 476 807
rect 477 803 479 807
rect 479 803 481 807
rect 482 803 483 807
rect 483 803 486 807
rect 976 903 977 907
rect 977 903 980 907
rect 981 903 983 907
rect 983 903 985 907
rect 986 903 987 907
rect 987 903 990 907
rect 472 603 473 607
rect 473 603 476 607
rect 477 603 479 607
rect 479 603 481 607
rect 482 603 483 607
rect 483 603 486 607
rect 894 528 898 532
rect 286 348 290 352
rect 78 258 82 262
rect 472 403 473 407
rect 473 403 476 407
rect 477 403 479 407
rect 479 403 481 407
rect 482 403 483 407
rect 483 403 486 407
rect 470 348 474 352
rect 454 258 458 262
rect 472 203 473 207
rect 473 203 476 207
rect 477 203 479 207
rect 479 203 481 207
rect 482 203 483 207
rect 483 203 486 207
rect 518 148 522 152
rect 558 258 562 262
rect 646 248 650 252
rect 718 148 722 152
rect 702 138 706 142
rect 878 138 882 142
rect 918 528 922 532
rect 1134 778 1138 782
rect 1142 778 1146 782
rect 976 703 977 707
rect 977 703 980 707
rect 981 703 983 707
rect 983 703 985 707
rect 986 703 987 707
rect 987 703 990 707
rect 976 503 977 507
rect 977 503 980 507
rect 981 503 983 507
rect 983 503 985 507
rect 986 503 987 507
rect 987 503 990 507
rect 918 448 922 452
rect 950 448 954 452
rect 1022 558 1026 562
rect 976 303 977 307
rect 977 303 980 307
rect 981 303 983 307
rect 983 303 985 307
rect 986 303 987 307
rect 987 303 990 307
rect 976 103 977 107
rect 977 103 980 107
rect 981 103 983 107
rect 983 103 985 107
rect 986 103 987 107
rect 987 103 990 107
rect 1134 558 1138 562
rect 472 3 473 7
rect 473 3 476 7
rect 477 3 479 7
rect 479 3 481 7
rect 482 3 483 7
rect 483 3 486 7
<< metal5 >>
rect 486 1203 488 1207
rect 472 1202 473 1203
rect 478 1202 480 1203
rect 485 1202 488 1203
rect 990 1103 992 1107
rect 976 1102 977 1103
rect 982 1102 984 1103
rect 989 1102 992 1103
rect 486 1003 488 1007
rect 472 1002 473 1003
rect 478 1002 480 1003
rect 485 1002 488 1003
rect 990 903 992 907
rect 976 902 977 903
rect 982 902 984 903
rect 989 902 992 903
rect 486 803 488 807
rect 472 802 473 803
rect 478 802 480 803
rect 485 802 488 803
rect 1138 778 1142 781
rect 990 703 992 707
rect 976 702 977 703
rect 982 702 984 703
rect 989 702 992 703
rect 486 603 488 607
rect 472 602 473 603
rect 478 602 480 603
rect 485 602 488 603
rect 1026 558 1134 561
rect 898 528 918 531
rect 990 503 992 507
rect 976 502 977 503
rect 982 502 984 503
rect 989 502 992 503
rect 922 448 950 451
rect 486 403 488 407
rect 472 402 473 403
rect 478 402 480 403
rect 485 402 488 403
rect 290 348 470 351
rect 990 303 992 307
rect 976 302 977 303
rect 982 302 984 303
rect 989 302 992 303
rect 82 258 454 261
rect 562 258 649 261
rect 646 252 649 258
rect 486 203 488 207
rect 472 202 473 203
rect 478 202 480 203
rect 485 202 488 203
rect 522 148 718 151
rect 706 138 878 141
rect 990 103 992 107
rect 976 102 977 103
rect 982 102 984 103
rect 989 102 992 103
rect 486 3 488 7
rect 472 2 473 3
rect 478 2 480 3
rect 485 2 488 3
<< m6contact >>
rect 473 1203 476 1207
rect 476 1203 477 1207
rect 477 1203 478 1207
rect 480 1203 481 1207
rect 481 1203 482 1207
rect 482 1203 485 1207
rect 473 1202 478 1203
rect 480 1202 485 1203
rect 977 1103 980 1107
rect 980 1103 981 1107
rect 981 1103 982 1107
rect 984 1103 985 1107
rect 985 1103 986 1107
rect 986 1103 989 1107
rect 977 1102 982 1103
rect 984 1102 989 1103
rect 473 1003 476 1007
rect 476 1003 477 1007
rect 477 1003 478 1007
rect 480 1003 481 1007
rect 481 1003 482 1007
rect 482 1003 485 1007
rect 473 1002 478 1003
rect 480 1002 485 1003
rect 977 903 980 907
rect 980 903 981 907
rect 981 903 982 907
rect 984 903 985 907
rect 985 903 986 907
rect 986 903 989 907
rect 977 902 982 903
rect 984 902 989 903
rect 473 803 476 807
rect 476 803 477 807
rect 477 803 478 807
rect 480 803 481 807
rect 481 803 482 807
rect 482 803 485 807
rect 473 802 478 803
rect 480 802 485 803
rect 977 703 980 707
rect 980 703 981 707
rect 981 703 982 707
rect 984 703 985 707
rect 985 703 986 707
rect 986 703 989 707
rect 977 702 982 703
rect 984 702 989 703
rect 473 603 476 607
rect 476 603 477 607
rect 477 603 478 607
rect 480 603 481 607
rect 481 603 482 607
rect 482 603 485 607
rect 473 602 478 603
rect 480 602 485 603
rect 977 503 980 507
rect 980 503 981 507
rect 981 503 982 507
rect 984 503 985 507
rect 985 503 986 507
rect 986 503 989 507
rect 977 502 982 503
rect 984 502 989 503
rect 473 403 476 407
rect 476 403 477 407
rect 477 403 478 407
rect 480 403 481 407
rect 481 403 482 407
rect 482 403 485 407
rect 473 402 478 403
rect 480 402 485 403
rect 977 303 980 307
rect 980 303 981 307
rect 981 303 982 307
rect 984 303 985 307
rect 985 303 986 307
rect 986 303 989 307
rect 977 302 982 303
rect 984 302 989 303
rect 473 203 476 207
rect 476 203 477 207
rect 477 203 478 207
rect 480 203 481 207
rect 481 203 482 207
rect 482 203 485 207
rect 473 202 478 203
rect 480 202 485 203
rect 977 103 980 107
rect 980 103 981 107
rect 981 103 982 107
rect 984 103 985 107
rect 985 103 986 107
rect 986 103 989 107
rect 977 102 982 103
rect 984 102 989 103
rect 473 3 476 7
rect 476 3 477 7
rect 477 3 478 7
rect 480 3 481 7
rect 481 3 482 7
rect 482 3 485 7
rect 473 2 478 3
rect 480 2 485 3
<< metal6 >>
rect 472 1207 488 1230
rect 472 1202 473 1207
rect 478 1202 480 1207
rect 485 1202 488 1207
rect 472 1007 488 1202
rect 472 1002 473 1007
rect 478 1002 480 1007
rect 485 1002 488 1007
rect 472 807 488 1002
rect 472 802 473 807
rect 478 802 480 807
rect 485 802 488 807
rect 472 607 488 802
rect 472 602 473 607
rect 478 602 480 607
rect 485 602 488 607
rect 472 407 488 602
rect 472 402 473 407
rect 478 402 480 407
rect 485 402 488 407
rect 472 207 488 402
rect 472 202 473 207
rect 478 202 480 207
rect 485 202 488 207
rect 472 7 488 202
rect 472 2 473 7
rect 478 2 480 7
rect 485 2 488 7
rect 472 -30 488 2
rect 976 1107 992 1230
rect 976 1102 977 1107
rect 982 1102 984 1107
rect 989 1102 992 1107
rect 976 907 992 1102
rect 976 902 977 907
rect 982 902 984 907
rect 989 902 992 907
rect 976 707 992 902
rect 976 702 977 707
rect 982 702 984 707
rect 989 702 992 707
rect 976 507 992 702
rect 976 502 977 507
rect 982 502 984 507
rect 989 502 992 507
rect 976 307 992 502
rect 976 302 977 307
rect 982 302 984 307
rect 989 302 992 307
rect 976 107 992 302
rect 976 102 977 107
rect 982 102 984 107
rect 989 102 992 107
rect 976 -30 992 102
use DFFPOSX1  DFFPOSX1_39
timestamp 1537603335
transform -1 0 100 0 1 1105
box 0 0 96 100
use BUFX2  BUFX2_12
timestamp 1537603335
transform -1 0 124 0 1 1105
box 0 0 24 100
use XNOR2X1  XNOR2X1_11
timestamp 1537603335
transform -1 0 180 0 1 1105
box 0 0 56 100
use INVX1  INVX1_27
timestamp 1537603335
transform 1 0 180 0 1 1105
box 0 0 16 100
use BUFX2  BUFX2_15
timestamp 1537603335
transform 1 0 196 0 1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_42
timestamp 1537603335
transform -1 0 316 0 1 1105
box 0 0 96 100
use XOR2X1  XOR2X1_5
timestamp 1537603335
transform -1 0 372 0 1 1105
box 0 0 56 100
use OAI21X1  OAI21X1_42
timestamp 1537603335
transform 1 0 372 0 1 1105
box 0 0 32 100
use AOI21X1  AOI21X1_21
timestamp 1537603335
transform 1 0 404 0 1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_41
timestamp 1537603335
transform -1 0 460 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_10
timestamp 1537603335
transform 1 0 460 0 1 1105
box 0 0 24 100
use FILL  FILL_11_0_0
timestamp 1537603335
transform -1 0 492 0 1 1105
box 0 0 8 100
use FILL  FILL_11_0_1
timestamp 1537603335
transform -1 0 500 0 1 1105
box 0 0 8 100
use NOR3X1  NOR3X1_8
timestamp 1537603335
transform -1 0 564 0 1 1105
box 0 0 64 100
use NOR2X1  NOR2X1_40
timestamp 1537603335
transform -1 0 588 0 1 1105
box 0 0 24 100
use XNOR2X1  XNOR2X1_12
timestamp 1537603335
transform 1 0 588 0 1 1105
box 0 0 56 100
use NAND2X1  NAND2X1_28
timestamp 1537603335
transform -1 0 668 0 1 1105
box 0 0 24 100
use INVX2  INVX2_9
timestamp 1537603335
transform -1 0 684 0 1 1105
box 0 0 16 100
use BUFX2  BUFX2_14
timestamp 1537603335
transform 1 0 684 0 1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_40
timestamp 1537603335
transform 1 0 708 0 1 1105
box 0 0 96 100
use BUFX2  BUFX2_13
timestamp 1537603335
transform 1 0 804 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_7
timestamp 1537603335
transform 1 0 828 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_49
timestamp 1537603335
transform 1 0 852 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_37
timestamp 1537603335
transform 1 0 876 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_39
timestamp 1537603335
transform 1 0 900 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_53
timestamp 1537603335
transform 1 0 924 0 1 1105
box 0 0 24 100
use XOR2X1  XOR2X1_2
timestamp 1537603335
transform 1 0 948 0 1 1105
box 0 0 56 100
use FILL  FILL_11_1_0
timestamp 1537603335
transform 1 0 1004 0 1 1105
box 0 0 8 100
use FILL  FILL_11_1_1
timestamp 1537603335
transform 1 0 1012 0 1 1105
box 0 0 8 100
use BUFX2  BUFX2_16
timestamp 1537603335
transform 1 0 1020 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_57
timestamp 1537603335
transform 1 0 1044 0 1 1105
box 0 0 24 100
use NAND2X1  NAND2X1_8
timestamp 1537603335
transform 1 0 1068 0 1 1105
box 0 0 24 100
use NAND2X1  NAND2X1_17
timestamp 1537603335
transform 1 0 1092 0 1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_3
timestamp 1537603335
transform 1 0 1116 0 1 1105
box 0 0 96 100
use BUFX2  BUFX2_18
timestamp 1537603335
transform 1 0 1212 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_19
timestamp 1537603335
transform -1 0 1260 0 1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_4
timestamp 1537603335
transform -1 0 1356 0 1 1105
box 0 0 96 100
use BUFX2  BUFX2_28
timestamp 1537603335
transform 1 0 1356 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_65
timestamp 1537603335
transform -1 0 1404 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_45
timestamp 1537603335
transform 1 0 1404 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_36
timestamp 1537603335
transform 1 0 1428 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_48
timestamp 1537603335
transform 1 0 1452 0 1 1105
box 0 0 24 100
use FILL  FILL_12_1
timestamp 1537603335
transform 1 0 1476 0 1 1105
box 0 0 8 100
use BUFX2  BUFX2_27
timestamp 1537603335
transform -1 0 28 0 -1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_12
timestamp 1537603335
transform -1 0 124 0 -1 1105
box 0 0 96 100
use INVX1  INVX1_15
timestamp 1537603335
transform 1 0 124 0 -1 1105
box 0 0 16 100
use NOR2X1  NOR2X1_27
timestamp 1537603335
transform 1 0 140 0 -1 1105
box 0 0 24 100
use BUFX2  BUFX2_11
timestamp 1537603335
transform -1 0 188 0 -1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_38
timestamp 1537603335
transform -1 0 284 0 -1 1105
box 0 0 96 100
use XNOR2X1  XNOR2X1_10
timestamp 1537603335
transform -1 0 340 0 -1 1105
box 0 0 56 100
use NOR3X1  NOR3X1_6
timestamp 1537603335
transform -1 0 404 0 -1 1105
box 0 0 64 100
use INVX1  INVX1_26
timestamp 1537603335
transform 1 0 404 0 -1 1105
box 0 0 16 100
use AND2X2  AND2X2_14
timestamp 1537603335
transform -1 0 452 0 -1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_41
timestamp 1537603335
transform -1 0 484 0 -1 1105
box 0 0 32 100
use FILL  FILL_10_0_0
timestamp 1537603335
transform 1 0 484 0 -1 1105
box 0 0 8 100
use FILL  FILL_10_0_1
timestamp 1537603335
transform 1 0 492 0 -1 1105
box 0 0 8 100
use NOR3X1  NOR3X1_7
timestamp 1537603335
transform 1 0 500 0 -1 1105
box 0 0 64 100
use OAI21X1  OAI21X1_45
timestamp 1537603335
transform -1 0 596 0 -1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_43
timestamp 1537603335
transform -1 0 628 0 -1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_30
timestamp 1537603335
transform -1 0 652 0 -1 1105
box 0 0 24 100
use NAND2X1  NAND2X1_29
timestamp 1537603335
transform 1 0 652 0 -1 1105
box 0 0 24 100
use XNOR2X1  XNOR2X1_13
timestamp 1537603335
transform 1 0 676 0 -1 1105
box 0 0 56 100
use INVX1  INVX1_28
timestamp 1537603335
transform -1 0 748 0 -1 1105
box 0 0 16 100
use DFFPOSX1  DFFPOSX1_41
timestamp 1537603335
transform -1 0 844 0 -1 1105
box 0 0 96 100
use BUFX2  BUFX2_31
timestamp 1537603335
transform 1 0 844 0 -1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_19
timestamp 1537603335
transform 1 0 868 0 -1 1105
box 0 0 96 100
use FILL  FILL_10_1_0
timestamp 1537603335
transform 1 0 964 0 -1 1105
box 0 0 8 100
use FILL  FILL_10_1_1
timestamp 1537603335
transform 1 0 972 0 -1 1105
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_26
timestamp 1537603335
transform 1 0 980 0 -1 1105
box 0 0 96 100
use INVX1  INVX1_5
timestamp 1537603335
transform 1 0 1076 0 -1 1105
box 0 0 16 100
use MUX2X1  MUX2X1_1
timestamp 1537603335
transform 1 0 1092 0 -1 1105
box 0 0 48 100
use OAI21X1  OAI21X1_3
timestamp 1537603335
transform -1 0 1172 0 -1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_3
timestamp 1537603335
transform 1 0 1172 0 -1 1105
box 0 0 48 100
use AOI21X1  AOI21X1_8
timestamp 1537603335
transform 1 0 1220 0 -1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_18
timestamp 1537603335
transform 1 0 1252 0 -1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_4
timestamp 1537603335
transform 1 0 1276 0 -1 1105
box 0 0 32 100
use AOI21X1  AOI21X1_9
timestamp 1537603335
transform 1 0 1308 0 -1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_19
timestamp 1537603335
transform 1 0 1340 0 -1 1105
box 0 0 24 100
use NOR2X1  NOR2X1_28
timestamp 1537603335
transform -1 0 1388 0 -1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_13
timestamp 1537603335
transform 1 0 1388 0 -1 1105
box 0 0 96 100
use BUFX2  BUFX2_2
timestamp 1537603335
transform -1 0 28 0 1 905
box 0 0 24 100
use BUFX2  BUFX2_3
timestamp 1537603335
transform -1 0 52 0 1 905
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_30
timestamp 1537603335
transform -1 0 148 0 1 905
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_29
timestamp 1537603335
transform -1 0 244 0 1 905
box 0 0 96 100
use XNOR2X1  XNOR2X1_2
timestamp 1537603335
transform -1 0 300 0 1 905
box 0 0 56 100
use OAI21X1  OAI21X1_31
timestamp 1537603335
transform 1 0 300 0 1 905
box 0 0 32 100
use NOR2X1  NOR2X1_34
timestamp 1537603335
transform 1 0 332 0 1 905
box 0 0 24 100
use XOR2X1  XOR2X1_4
timestamp 1537603335
transform -1 0 412 0 1 905
box 0 0 56 100
use NOR2X1  NOR2X1_39
timestamp 1537603335
transform -1 0 436 0 1 905
box 0 0 24 100
use OAI21X1  OAI21X1_40
timestamp 1537603335
transform 1 0 436 0 1 905
box 0 0 32 100
use FILL  FILL_9_0_0
timestamp 1537603335
transform -1 0 476 0 1 905
box 0 0 8 100
use FILL  FILL_9_0_1
timestamp 1537603335
transform -1 0 484 0 1 905
box 0 0 8 100
use AOI21X1  AOI21X1_20
timestamp 1537603335
transform -1 0 516 0 1 905
box 0 0 32 100
use AOI21X1  AOI21X1_19
timestamp 1537603335
transform -1 0 548 0 1 905
box 0 0 32 100
use INVX1  INVX1_29
timestamp 1537603335
transform -1 0 564 0 1 905
box 0 0 16 100
use NAND3X1  NAND3X1_14
timestamp 1537603335
transform 1 0 564 0 1 905
box 0 0 32 100
use BUFX2  BUFX2_8
timestamp 1537603335
transform 1 0 596 0 1 905
box 0 0 24 100
use AOI21X1  AOI21X1_22
timestamp 1537603335
transform 1 0 620 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_44
timestamp 1537603335
transform -1 0 684 0 1 905
box 0 0 32 100
use INVX1  INVX1_19
timestamp 1537603335
transform 1 0 684 0 1 905
box 0 0 16 100
use NOR2X1  NOR2X1_31
timestamp 1537603335
transform 1 0 700 0 1 905
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_16
timestamp 1537603335
transform 1 0 724 0 1 905
box 0 0 96 100
use BUFX2  BUFX2_61
timestamp 1537603335
transform 1 0 820 0 1 905
box 0 0 24 100
use BUFX2  BUFX2_70
timestamp 1537603335
transform -1 0 868 0 1 905
box 0 0 24 100
use MUX2X1  MUX2X1_2
timestamp 1537603335
transform -1 0 916 0 1 905
box 0 0 48 100
use BUFX2  BUFX2_71
timestamp 1537603335
transform 1 0 916 0 1 905
box 0 0 24 100
use NOR2X1  NOR2X1_13
timestamp 1537603335
transform 1 0 940 0 1 905
box 0 0 24 100
use INVX2  INVX2_4
timestamp 1537603335
transform -1 0 980 0 1 905
box 0 0 16 100
use FILL  FILL_9_1_0
timestamp 1537603335
transform -1 0 988 0 1 905
box 0 0 8 100
use FILL  FILL_9_1_1
timestamp 1537603335
transform -1 0 996 0 1 905
box 0 0 8 100
use BUFX2  BUFX2_54
timestamp 1537603335
transform -1 0 1020 0 1 905
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_20
timestamp 1537603335
transform -1 0 1116 0 1 905
box 0 0 96 100
use OAI21X1  OAI21X1_22
timestamp 1537603335
transform -1 0 1148 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_21
timestamp 1537603335
transform -1 0 1180 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_9
timestamp 1537603335
transform 1 0 1180 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_24
timestamp 1537603335
transform 1 0 1212 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_23
timestamp 1537603335
transform 1 0 1244 0 1 905
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_24
timestamp 1537603335
transform 1 0 1276 0 1 905
box 0 0 96 100
use AOI21X1  AOI21X1_4
timestamp 1537603335
transform -1 0 1404 0 1 905
box 0 0 32 100
use BUFX2  BUFX2_58
timestamp 1537603335
transform 1 0 1404 0 1 905
box 0 0 24 100
use INVX1  INVX1_11
timestamp 1537603335
transform -1 0 1444 0 1 905
box 0 0 16 100
use BUFX2  BUFX2_44
timestamp 1537603335
transform 1 0 1444 0 1 905
box 0 0 24 100
use FILL  FILL_10_1
timestamp 1537603335
transform 1 0 1468 0 1 905
box 0 0 8 100
use FILL  FILL_10_2
timestamp 1537603335
transform 1 0 1476 0 1 905
box 0 0 8 100
use BUFX2  BUFX2_9
timestamp 1537603335
transform -1 0 28 0 -1 905
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_36
timestamp 1537603335
transform -1 0 124 0 -1 905
box 0 0 96 100
use XNOR2X1  XNOR2X1_3
timestamp 1537603335
transform -1 0 180 0 -1 905
box 0 0 56 100
use OAI21X1  OAI21X1_32
timestamp 1537603335
transform 1 0 180 0 -1 905
box 0 0 32 100
use BUFX4  BUFX4_9
timestamp 1537603335
transform 1 0 212 0 -1 905
box 0 0 32 100
use INVX1  INVX1_21
timestamp 1537603335
transform 1 0 244 0 -1 905
box 0 0 16 100
use NOR2X1  NOR2X1_33
timestamp 1537603335
transform -1 0 284 0 -1 905
box 0 0 24 100
use XNOR2X1  XNOR2X1_9
timestamp 1537603335
transform -1 0 340 0 -1 905
box 0 0 56 100
use DFFPOSX1  DFFPOSX1_37
timestamp 1537603335
transform 1 0 340 0 -1 905
box 0 0 96 100
use NAND3X1  NAND3X1_13
timestamp 1537603335
transform -1 0 468 0 -1 905
box 0 0 32 100
use FILL  FILL_8_0_0
timestamp 1537603335
transform -1 0 476 0 -1 905
box 0 0 8 100
use FILL  FILL_8_0_1
timestamp 1537603335
transform -1 0 484 0 -1 905
box 0 0 8 100
use OAI21X1  OAI21X1_38
timestamp 1537603335
transform -1 0 516 0 -1 905
box 0 0 32 100
use OAI21X1  OAI21X1_39
timestamp 1537603335
transform -1 0 548 0 -1 905
box 0 0 32 100
use INVX2  INVX2_8
timestamp 1537603335
transform -1 0 564 0 -1 905
box 0 0 16 100
use INVX1  INVX1_25
timestamp 1537603335
transform 1 0 564 0 -1 905
box 0 0 16 100
use NAND3X1  NAND3X1_12
timestamp 1537603335
transform -1 0 612 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_13
timestamp 1537603335
transform -1 0 644 0 -1 905
box 0 0 32 100
use INVX1  INVX1_24
timestamp 1537603335
transform -1 0 660 0 -1 905
box 0 0 16 100
use OAI21X1  OAI21X1_37
timestamp 1537603335
transform 1 0 660 0 -1 905
box 0 0 32 100
use BUFX4  BUFX4_5
timestamp 1537603335
transform -1 0 724 0 -1 905
box 0 0 32 100
use XNOR2X1  XNOR2X1_8
timestamp 1537603335
transform 1 0 724 0 -1 905
box 0 0 56 100
use DFFPOSX1  DFFPOSX1_35
timestamp 1537603335
transform -1 0 876 0 -1 905
box 0 0 96 100
use BUFX4  BUFX4_19
timestamp 1537603335
transform 1 0 876 0 -1 905
box 0 0 32 100
use BUFX2  BUFX2_74
timestamp 1537603335
transform 1 0 908 0 -1 905
box 0 0 24 100
use BUFX4  BUFX4_12
timestamp 1537603335
transform 1 0 932 0 -1 905
box 0 0 32 100
use OAI21X1  OAI21X1_20
timestamp 1537603335
transform -1 0 996 0 -1 905
box 0 0 32 100
use FILL  FILL_8_1_0
timestamp 1537603335
transform 1 0 996 0 -1 905
box 0 0 8 100
use FILL  FILL_8_1_1
timestamp 1537603335
transform 1 0 1004 0 -1 905
box 0 0 8 100
use BUFX4  BUFX4_11
timestamp 1537603335
transform 1 0 1012 0 -1 905
box 0 0 32 100
use INVX4  INVX4_1
timestamp 1537603335
transform 1 0 1044 0 -1 905
box 0 0 24 100
use OAI21X1  OAI21X1_5
timestamp 1537603335
transform 1 0 1068 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_3
timestamp 1537603335
transform 1 0 1100 0 -1 905
box 0 0 32 100
use OAI22X1  OAI22X1_1
timestamp 1537603335
transform -1 0 1172 0 -1 905
box 0 0 40 100
use NAND3X1  NAND3X1_7
timestamp 1537603335
transform -1 0 1204 0 -1 905
box 0 0 32 100
use INVX4  INVX4_2
timestamp 1537603335
transform 1 0 1204 0 -1 905
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_23
timestamp 1537603335
transform -1 0 1324 0 -1 905
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_25
timestamp 1537603335
transform 1 0 1324 0 -1 905
box 0 0 96 100
use BUFX4  BUFX4_18
timestamp 1537603335
transform -1 0 1452 0 -1 905
box 0 0 32 100
use BUFX2  BUFX2_59
timestamp 1537603335
transform 1 0 1452 0 -1 905
box 0 0 24 100
use FILL  FILL_9_1
timestamp 1537603335
transform -1 0 1484 0 -1 905
box 0 0 8 100
use BUFX2  BUFX2_1
timestamp 1537603335
transform -1 0 28 0 1 705
box 0 0 24 100
use NOR3X1  NOR3X1_4
timestamp 1537603335
transform -1 0 92 0 1 705
box 0 0 64 100
use AND2X2  AND2X2_12
timestamp 1537603335
transform 1 0 92 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_11
timestamp 1537603335
transform 1 0 124 0 1 705
box 0 0 32 100
use NAND2X1  NAND2X1_20
timestamp 1537603335
transform 1 0 156 0 1 705
box 0 0 24 100
use NAND3X1  NAND3X1_9
timestamp 1537603335
transform -1 0 212 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_2
timestamp 1537603335
transform -1 0 244 0 1 705
box 0 0 32 100
use NAND2X1  NAND2X1_21
timestamp 1537603335
transform 1 0 244 0 1 705
box 0 0 24 100
use BUFX4  BUFX4_6
timestamp 1537603335
transform -1 0 300 0 1 705
box 0 0 32 100
use NOR2X1  NOR2X1_37
timestamp 1537603335
transform 1 0 300 0 1 705
box 0 0 24 100
use NOR2X1  NOR2X1_36
timestamp 1537603335
transform 1 0 324 0 1 705
box 0 0 24 100
use OR2X2  OR2X2_3
timestamp 1537603335
transform -1 0 380 0 1 705
box 0 0 32 100
use NOR2X1  NOR2X1_35
timestamp 1537603335
transform -1 0 404 0 1 705
box 0 0 24 100
use NAND2X1  NAND2X1_27
timestamp 1537603335
transform -1 0 428 0 1 705
box 0 0 24 100
use NOR2X1  NOR2X1_38
timestamp 1537603335
transform -1 0 452 0 1 705
box 0 0 24 100
use NAND2X1  NAND2X1_26
timestamp 1537603335
transform 1 0 452 0 1 705
box 0 0 24 100
use FILL  FILL_7_0_0
timestamp 1537603335
transform 1 0 476 0 1 705
box 0 0 8 100
use FILL  FILL_7_0_1
timestamp 1537603335
transform 1 0 484 0 1 705
box 0 0 8 100
use INVX1  INVX1_23
timestamp 1537603335
transform 1 0 492 0 1 705
box 0 0 16 100
use AOI21X1  AOI21X1_18
timestamp 1537603335
transform 1 0 508 0 1 705
box 0 0 32 100
use AOI21X1  AOI21X1_17
timestamp 1537603335
transform -1 0 572 0 1 705
box 0 0 32 100
use INVX8  INVX8_1
timestamp 1537603335
transform 1 0 572 0 1 705
box 0 0 40 100
use DFFPOSX1  DFFPOSX1_34
timestamp 1537603335
transform -1 0 708 0 1 705
box 0 0 96 100
use XNOR2X1  XNOR2X1_1
timestamp 1537603335
transform -1 0 764 0 1 705
box 0 0 56 100
use NOR2X1  NOR2X1_14
timestamp 1537603335
transform -1 0 788 0 1 705
box 0 0 24 100
use NAND2X1  NAND2X1_11
timestamp 1537603335
transform 1 0 788 0 1 705
box 0 0 24 100
use AND2X2  AND2X2_6
timestamp 1537603335
transform -1 0 844 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_6
timestamp 1537603335
transform 1 0 844 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_4
timestamp 1537603335
transform -1 0 908 0 1 705
box 0 0 32 100
use MUX2X1  MUX2X1_4
timestamp 1537603335
transform 1 0 908 0 1 705
box 0 0 48 100
use NAND3X1  NAND3X1_5
timestamp 1537603335
transform 1 0 956 0 1 705
box 0 0 32 100
use FILL  FILL_7_1_0
timestamp 1537603335
transform -1 0 996 0 1 705
box 0 0 8 100
use FILL  FILL_7_1_1
timestamp 1537603335
transform -1 0 1004 0 1 705
box 0 0 8 100
use NOR3X1  NOR3X1_2
timestamp 1537603335
transform -1 0 1068 0 1 705
box 0 0 64 100
use NAND3X1  NAND3X1_8
timestamp 1537603335
transform -1 0 1100 0 1 705
box 0 0 32 100
use OAI21X1  OAI21X1_25
timestamp 1537603335
transform 1 0 1100 0 1 705
box 0 0 32 100
use OAI21X1  OAI21X1_15
timestamp 1537603335
transform 1 0 1132 0 1 705
box 0 0 32 100
use AOI21X1  AOI21X1_5
timestamp 1537603335
transform -1 0 1196 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_10
timestamp 1537603335
transform 1 0 1196 0 1 705
box 0 0 32 100
use OAI21X1  OAI21X1_16
timestamp 1537603335
transform 1 0 1228 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_7
timestamp 1537603335
transform 1 0 1260 0 1 705
box 0 0 32 100
use OAI21X1  OAI21X1_19
timestamp 1537603335
transform 1 0 1292 0 1 705
box 0 0 32 100
use INVX2  INVX2_2
timestamp 1537603335
transform 1 0 1324 0 1 705
box 0 0 16 100
use OAI21X1  OAI21X1_17
timestamp 1537603335
transform 1 0 1340 0 1 705
box 0 0 32 100
use OAI21X1  OAI21X1_18
timestamp 1537603335
transform 1 0 1372 0 1 705
box 0 0 32 100
use AOI21X1  AOI21X1_3
timestamp 1537603335
transform -1 0 1436 0 1 705
box 0 0 32 100
use BUFX2  BUFX2_56
timestamp 1537603335
transform 1 0 1436 0 1 705
box 0 0 24 100
use FILL  FILL_8_1
timestamp 1537603335
transform 1 0 1460 0 1 705
box 0 0 8 100
use FILL  FILL_8_2
timestamp 1537603335
transform 1 0 1468 0 1 705
box 0 0 8 100
use FILL  FILL_8_3
timestamp 1537603335
transform 1 0 1476 0 1 705
box 0 0 8 100
use BUFX2  BUFX2_4
timestamp 1537603335
transform -1 0 28 0 -1 705
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_31
timestamp 1537603335
transform -1 0 124 0 -1 705
box 0 0 96 100
use INVX2  INVX2_7
timestamp 1537603335
transform 1 0 124 0 -1 705
box 0 0 16 100
use XNOR2X1  XNOR2X1_4
timestamp 1537603335
transform -1 0 196 0 -1 705
box 0 0 56 100
use AOI21X1  AOI21X1_15
timestamp 1537603335
transform 1 0 196 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_33
timestamp 1537603335
transform -1 0 260 0 -1 705
box 0 0 32 100
use NAND3X1  NAND3X1_10
timestamp 1537603335
transform -1 0 292 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_34
timestamp 1537603335
transform -1 0 324 0 -1 705
box 0 0 32 100
use NAND3X1  NAND3X1_11
timestamp 1537603335
transform 1 0 324 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_35
timestamp 1537603335
transform -1 0 388 0 -1 705
box 0 0 32 100
use INVX1  INVX1_22
timestamp 1537603335
transform -1 0 404 0 -1 705
box 0 0 16 100
use NAND2X1  NAND2X1_24
timestamp 1537603335
transform -1 0 428 0 -1 705
box 0 0 24 100
use NAND2X1  NAND2X1_23
timestamp 1537603335
transform 1 0 428 0 -1 705
box 0 0 24 100
use AOI21X1  AOI21X1_16
timestamp 1537603335
transform -1 0 484 0 -1 705
box 0 0 32 100
use FILL  FILL_6_0_0
timestamp 1537603335
transform -1 0 492 0 -1 705
box 0 0 8 100
use FILL  FILL_6_0_1
timestamp 1537603335
transform -1 0 500 0 -1 705
box 0 0 8 100
use NOR3X1  NOR3X1_5
timestamp 1537603335
transform -1 0 564 0 -1 705
box 0 0 64 100
use OAI21X1  OAI21X1_36
timestamp 1537603335
transform 1 0 564 0 -1 705
box 0 0 32 100
use NAND2X1  NAND2X1_25
timestamp 1537603335
transform 1 0 596 0 -1 705
box 0 0 24 100
use BUFX4  BUFX4_2
timestamp 1537603335
transform -1 0 652 0 -1 705
box 0 0 32 100
use XNOR2X1  XNOR2X1_7
timestamp 1537603335
transform 1 0 652 0 -1 705
box 0 0 56 100
use BUFX4  BUFX4_4
timestamp 1537603335
transform 1 0 708 0 -1 705
box 0 0 32 100
use NOR3X1  NOR3X1_1
timestamp 1537603335
transform -1 0 804 0 -1 705
box 0 0 64 100
use NOR2X1  NOR2X1_9
timestamp 1537603335
transform -1 0 828 0 -1 705
box 0 0 24 100
use AND2X2  AND2X2_2
timestamp 1537603335
transform -1 0 860 0 -1 705
box 0 0 32 100
use NAND2X1  NAND2X1_14
timestamp 1537603335
transform 1 0 860 0 -1 705
box 0 0 24 100
use NAND2X1  NAND2X1_13
timestamp 1537603335
transform 1 0 884 0 -1 705
box 0 0 24 100
use NOR2X1  NOR2X1_15
timestamp 1537603335
transform 1 0 908 0 -1 705
box 0 0 24 100
use NOR3X1  NOR3X1_3
timestamp 1537603335
transform 1 0 932 0 -1 705
box 0 0 64 100
use FILL  FILL_6_1_0
timestamp 1537603335
transform -1 0 1004 0 -1 705
box 0 0 8 100
use FILL  FILL_6_1_1
timestamp 1537603335
transform -1 0 1012 0 -1 705
box 0 0 8 100
use AND2X2  AND2X2_8
timestamp 1537603335
transform -1 0 1044 0 -1 705
box 0 0 32 100
use NAND2X1  NAND2X1_18
timestamp 1537603335
transform -1 0 1068 0 -1 705
box 0 0 24 100
use NAND3X1  NAND3X1_2
timestamp 1537603335
transform -1 0 1100 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_26
timestamp 1537603335
transform 1 0 1100 0 -1 705
box 0 0 32 100
use NAND3X1  NAND3X1_3
timestamp 1537603335
transform -1 0 1164 0 -1 705
box 0 0 32 100
use NOR2X1  NOR2X1_8
timestamp 1537603335
transform 1 0 1164 0 -1 705
box 0 0 24 100
use NAND3X1  NAND3X1_1
timestamp 1537603335
transform 1 0 1188 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_27
timestamp 1537603335
transform 1 0 1220 0 -1 705
box 0 0 32 100
use INVX2  INVX2_1
timestamp 1537603335
transform -1 0 1268 0 -1 705
box 0 0 16 100
use OAI21X1  OAI21X1_30
timestamp 1537603335
transform 1 0 1268 0 -1 705
box 0 0 32 100
use AOI21X1  AOI21X1_2
timestamp 1537603335
transform -1 0 1332 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_29
timestamp 1537603335
transform -1 0 1364 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_28
timestamp 1537603335
transform 1 0 1364 0 -1 705
box 0 0 32 100
use INVX1  INVX1_9
timestamp 1537603335
transform -1 0 1412 0 -1 705
box 0 0 16 100
use NAND2X1  NAND2X1_19
timestamp 1537603335
transform 1 0 1412 0 -1 705
box 0 0 24 100
use INVX1  INVX1_7
timestamp 1537603335
transform -1 0 1452 0 -1 705
box 0 0 16 100
use BUFX2  BUFX2_47
timestamp 1537603335
transform 1 0 1452 0 -1 705
box 0 0 24 100
use FILL  FILL_7_1
timestamp 1537603335
transform -1 0 1484 0 -1 705
box 0 0 8 100
use BUFX2  BUFX2_29
timestamp 1537603335
transform -1 0 28 0 1 505
box 0 0 24 100
use BUFX2  BUFX2_35
timestamp 1537603335
transform -1 0 52 0 1 505
box 0 0 24 100
use INVX1  INVX1_17
timestamp 1537603335
transform 1 0 52 0 1 505
box 0 0 16 100
use BUFX2  BUFX2_63
timestamp 1537603335
transform -1 0 92 0 1 505
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_28
timestamp 1537603335
transform -1 0 188 0 1 505
box 0 0 96 100
use XOR2X1  XOR2X1_3
timestamp 1537603335
transform 1 0 188 0 1 505
box 0 0 56 100
use DFFPOSX1  DFFPOSX1_43
timestamp 1537603335
transform 1 0 244 0 1 505
box 0 0 96 100
use BUFX2  BUFX2_69
timestamp 1537603335
transform 1 0 340 0 1 505
box 0 0 24 100
use BUFX4  BUFX4_20
timestamp 1537603335
transform -1 0 396 0 1 505
box 0 0 32 100
use NAND2X1  NAND2X1_22
timestamp 1537603335
transform -1 0 420 0 1 505
box 0 0 24 100
use XNOR2X1  XNOR2X1_6
timestamp 1537603335
transform -1 0 476 0 1 505
box 0 0 56 100
use FILL  FILL_5_0_0
timestamp 1537603335
transform 1 0 476 0 1 505
box 0 0 8 100
use FILL  FILL_5_0_1
timestamp 1537603335
transform 1 0 484 0 1 505
box 0 0 8 100
use XNOR2X1  XNOR2X1_5
timestamp 1537603335
transform 1 0 492 0 1 505
box 0 0 56 100
use BUFX4  BUFX4_1
timestamp 1537603335
transform 1 0 548 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_1
timestamp 1537603335
transform -1 0 612 0 1 505
box 0 0 32 100
use NOR2X1  NOR2X1_3
timestamp 1537603335
transform 1 0 612 0 1 505
box 0 0 24 100
use INVX1  INVX1_2
timestamp 1537603335
transform -1 0 652 0 1 505
box 0 0 16 100
use NAND2X1  NAND2X1_2
timestamp 1537603335
transform -1 0 676 0 1 505
box 0 0 24 100
use BUFX4  BUFX4_3
timestamp 1537603335
transform -1 0 708 0 1 505
box 0 0 32 100
use NAND2X1  NAND2X1_3
timestamp 1537603335
transform 1 0 708 0 1 505
box 0 0 24 100
use NOR2X1  NOR2X1_4
timestamp 1537603335
transform 1 0 732 0 1 505
box 0 0 24 100
use NOR2X1  NOR2X1_2
timestamp 1537603335
transform -1 0 780 0 1 505
box 0 0 24 100
use BUFX4  BUFX4_17
timestamp 1537603335
transform -1 0 812 0 1 505
box 0 0 32 100
use OAI21X1  OAI21X1_6
timestamp 1537603335
transform 1 0 812 0 1 505
box 0 0 32 100
use NAND2X1  NAND2X1_10
timestamp 1537603335
transform -1 0 868 0 1 505
box 0 0 24 100
use INVX1  INVX1_8
timestamp 1537603335
transform 1 0 868 0 1 505
box 0 0 16 100
use NOR2X1  NOR2X1_16
timestamp 1537603335
transform -1 0 908 0 1 505
box 0 0 24 100
use AOI22X1  AOI22X1_2
timestamp 1537603335
transform -1 0 948 0 1 505
box 0 0 40 100
use FILL  FILL_5_1_0
timestamp 1537603335
transform -1 0 956 0 1 505
box 0 0 8 100
use FILL  FILL_5_1_1
timestamp 1537603335
transform -1 0 964 0 1 505
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_22
timestamp 1537603335
transform -1 0 1060 0 1 505
box 0 0 96 100
use NOR2X1  NOR2X1_10
timestamp 1537603335
transform -1 0 1084 0 1 505
box 0 0 24 100
use BUFX4  BUFX4_14
timestamp 1537603335
transform 1 0 1084 0 1 505
box 0 0 32 100
use OAI21X1  OAI21X1_11
timestamp 1537603335
transform -1 0 1148 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_5
timestamp 1537603335
transform 1 0 1148 0 1 505
box 0 0 32 100
use OAI21X1  OAI21X1_14
timestamp 1537603335
transform 1 0 1180 0 1 505
box 0 0 32 100
use OAI21X1  OAI21X1_13
timestamp 1537603335
transform -1 0 1244 0 1 505
box 0 0 32 100
use OAI21X1  OAI21X1_12
timestamp 1537603335
transform 1 0 1244 0 1 505
box 0 0 32 100
use NAND2X1  NAND2X1_15
timestamp 1537603335
transform 1 0 1276 0 1 505
box 0 0 24 100
use AOI21X1  AOI21X1_1
timestamp 1537603335
transform 1 0 1300 0 1 505
box 0 0 32 100
use AOI21X1  AOI21X1_6
timestamp 1537603335
transform -1 0 1364 0 1 505
box 0 0 32 100
use INVX1  INVX1_12
timestamp 1537603335
transform -1 0 1380 0 1 505
box 0 0 16 100
use BUFX2  BUFX2_55
timestamp 1537603335
transform 1 0 1380 0 1 505
box 0 0 24 100
use NAND2X1  NAND2X1_12
timestamp 1537603335
transform 1 0 1404 0 1 505
box 0 0 24 100
use BUFX2  BUFX2_22
timestamp 1537603335
transform 1 0 1428 0 1 505
box 0 0 24 100
use NAND2X1  NAND2X1_9
timestamp 1537603335
transform 1 0 1452 0 1 505
box 0 0 24 100
use FILL  FILL_6_1
timestamp 1537603335
transform 1 0 1476 0 1 505
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_14
timestamp 1537603335
transform -1 0 100 0 -1 505
box 0 0 96 100
use NOR2X1  NOR2X1_29
timestamp 1537603335
transform 1 0 100 0 -1 505
box 0 0 24 100
use BUFX2  BUFX2_75
timestamp 1537603335
transform 1 0 124 0 -1 505
box 0 0 24 100
use BUFX2  BUFX2_64
timestamp 1537603335
transform -1 0 172 0 -1 505
box 0 0 24 100
use BUFX4  BUFX4_8
timestamp 1537603335
transform -1 0 204 0 -1 505
box 0 0 32 100
use BUFX2  BUFX2_73
timestamp 1537603335
transform 1 0 204 0 -1 505
box 0 0 24 100
use INVX4  INVX4_3
timestamp 1537603335
transform -1 0 252 0 -1 505
box 0 0 24 100
use INVX1  INVX1_32
timestamp 1537603335
transform 1 0 252 0 -1 505
box 0 0 16 100
use NAND3X1  NAND3X1_19
timestamp 1537603335
transform -1 0 300 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_16
timestamp 1537603335
transform 1 0 300 0 -1 505
box 0 0 32 100
use NAND3X1  NAND3X1_17
timestamp 1537603335
transform 1 0 332 0 -1 505
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_33
timestamp 1537603335
transform -1 0 460 0 -1 505
box 0 0 96 100
use FILL  FILL_4_0_0
timestamp 1537603335
transform 1 0 460 0 -1 505
box 0 0 8 100
use FILL  FILL_4_0_1
timestamp 1537603335
transform 1 0 468 0 -1 505
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_32
timestamp 1537603335
transform 1 0 476 0 -1 505
box 0 0 96 100
use BUFX2  BUFX2_6
timestamp 1537603335
transform 1 0 572 0 -1 505
box 0 0 24 100
use BUFX2  BUFX2_5
timestamp 1537603335
transform 1 0 596 0 -1 505
box 0 0 24 100
use INVX1  INVX1_3
timestamp 1537603335
transform 1 0 620 0 -1 505
box 0 0 16 100
use NAND2X1  NAND2X1_5
timestamp 1537603335
transform -1 0 660 0 -1 505
box 0 0 24 100
use OR2X2  OR2X2_1
timestamp 1537603335
transform 1 0 660 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_1
timestamp 1537603335
transform 1 0 692 0 -1 505
box 0 0 24 100
use INVX1  INVX1_1
timestamp 1537603335
transform -1 0 732 0 -1 505
box 0 0 16 100
use NOR2X1  NOR2X1_7
timestamp 1537603335
transform 1 0 732 0 -1 505
box 0 0 24 100
use NOR2X1  NOR2X1_1
timestamp 1537603335
transform -1 0 780 0 -1 505
box 0 0 24 100
use NAND2X1  NAND2X1_6
timestamp 1537603335
transform 1 0 780 0 -1 505
box 0 0 24 100
use INVX2  INVX2_3
timestamp 1537603335
transform -1 0 820 0 -1 505
box 0 0 16 100
use NOR2X1  NOR2X1_12
timestamp 1537603335
transform 1 0 820 0 -1 505
box 0 0 24 100
use NAND2X1  NAND2X1_7
timestamp 1537603335
transform -1 0 868 0 -1 505
box 0 0 24 100
use OAI21X1  OAI21X1_1
timestamp 1537603335
transform -1 0 900 0 -1 505
box 0 0 32 100
use AOI22X1  AOI22X1_1
timestamp 1537603335
transform 1 0 900 0 -1 505
box 0 0 40 100
use OAI21X1  OAI21X1_2
timestamp 1537603335
transform -1 0 972 0 -1 505
box 0 0 32 100
use INVX1  INVX1_4
timestamp 1537603335
transform -1 0 988 0 -1 505
box 0 0 16 100
use FILL  FILL_4_1_0
timestamp 1537603335
transform -1 0 996 0 -1 505
box 0 0 8 100
use FILL  FILL_4_1_1
timestamp 1537603335
transform -1 0 1004 0 -1 505
box 0 0 8 100
use NOR2X1  NOR2X1_11
timestamp 1537603335
transform -1 0 1028 0 -1 505
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_18
timestamp 1537603335
transform -1 0 1124 0 -1 505
box 0 0 96 100
use INVX2  INVX2_6
timestamp 1537603335
transform 1 0 1124 0 -1 505
box 0 0 16 100
use BUFX4  BUFX4_15
timestamp 1537603335
transform 1 0 1140 0 -1 505
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_6
timestamp 1537603335
transform 1 0 1172 0 -1 505
box 0 0 96 100
use AOI21X1  AOI21X1_11
timestamp 1537603335
transform 1 0 1268 0 -1 505
box 0 0 32 100
use NOR2X1  NOR2X1_21
timestamp 1537603335
transform 1 0 1300 0 -1 505
box 0 0 24 100
use OAI21X1  OAI21X1_9
timestamp 1537603335
transform -1 0 1356 0 -1 505
box 0 0 32 100
use INVX1  INVX1_6
timestamp 1537603335
transform 1 0 1356 0 -1 505
box 0 0 16 100
use OAI21X1  OAI21X1_8
timestamp 1537603335
transform 1 0 1372 0 -1 505
box 0 0 32 100
use BUFX2  BUFX2_21
timestamp 1537603335
transform 1 0 1404 0 -1 505
box 0 0 24 100
use BUFX2  BUFX2_62
timestamp 1537603335
transform -1 0 1452 0 -1 505
box 0 0 24 100
use INVX1  INVX1_10
timestamp 1537603335
transform -1 0 1468 0 -1 505
box 0 0 16 100
use FILL  FILL_5_1
timestamp 1537603335
transform -1 0 1476 0 -1 505
box 0 0 8 100
use FILL  FILL_5_2
timestamp 1537603335
transform -1 0 1484 0 -1 505
box 0 0 8 100
use BUFX2  BUFX2_25
timestamp 1537603335
transform -1 0 28 0 1 305
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_10
timestamp 1537603335
transform -1 0 124 0 1 305
box 0 0 96 100
use INVX1  INVX1_13
timestamp 1537603335
transform 1 0 124 0 1 305
box 0 0 16 100
use NOR2X1  NOR2X1_25
timestamp 1537603335
transform 1 0 140 0 1 305
box 0 0 24 100
use NAND2X1  NAND2X1_37
timestamp 1537603335
transform 1 0 164 0 1 305
box 0 0 24 100
use NAND2X1  NAND2X1_32
timestamp 1537603335
transform -1 0 212 0 1 305
box 0 0 24 100
use NAND3X1  NAND3X1_20
timestamp 1537603335
transform -1 0 244 0 1 305
box 0 0 32 100
use NOR3X1  NOR3X1_12
timestamp 1537603335
transform -1 0 308 0 1 305
box 0 0 64 100
use NOR2X1  NOR2X1_49
timestamp 1537603335
transform 1 0 308 0 1 305
box 0 0 24 100
use NOR2X1  NOR2X1_51
timestamp 1537603335
transform -1 0 356 0 1 305
box 0 0 24 100
use INVX1  INVX1_34
timestamp 1537603335
transform -1 0 372 0 1 305
box 0 0 16 100
use OAI21X1  OAI21X1_58
timestamp 1537603335
transform 1 0 372 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_4
timestamp 1537603335
transform -1 0 436 0 1 305
box 0 0 32 100
use NAND2X1  NAND2X1_34
timestamp 1537603335
transform 1 0 436 0 1 305
box 0 0 24 100
use INVX1  INVX1_37
timestamp 1537603335
transform 1 0 460 0 1 305
box 0 0 16 100
use FILL  FILL_3_0_0
timestamp 1537603335
transform -1 0 484 0 1 305
box 0 0 8 100
use FILL  FILL_3_0_1
timestamp 1537603335
transform -1 0 492 0 1 305
box 0 0 8 100
use OAI21X1  OAI21X1_59
timestamp 1537603335
transform -1 0 524 0 1 305
box 0 0 32 100
use OAI21X1  OAI21X1_49
timestamp 1537603335
transform -1 0 556 0 1 305
box 0 0 32 100
use NOR2X1  NOR2X1_50
timestamp 1537603335
transform 1 0 556 0 1 305
box 0 0 24 100
use OAI21X1  OAI21X1_50
timestamp 1537603335
transform -1 0 612 0 1 305
box 0 0 32 100
use INVX4  INVX4_4
timestamp 1537603335
transform -1 0 636 0 1 305
box 0 0 24 100
use NAND2X1  NAND2X1_36
timestamp 1537603335
transform 1 0 636 0 1 305
box 0 0 24 100
use NOR3X1  NOR3X1_14
timestamp 1537603335
transform 1 0 660 0 1 305
box 0 0 64 100
use NAND2X1  NAND2X1_38
timestamp 1537603335
transform -1 0 748 0 1 305
box 0 0 24 100
use NAND3X1  NAND3X1_18
timestamp 1537603335
transform 1 0 748 0 1 305
box 0 0 32 100
use INVX1  INVX1_36
timestamp 1537603335
transform 1 0 780 0 1 305
box 0 0 16 100
use AOI21X1  AOI21X1_26
timestamp 1537603335
transform 1 0 796 0 1 305
box 0 0 32 100
use NOR2X1  NOR2X1_59
timestamp 1537603335
transform 1 0 828 0 1 305
box 0 0 24 100
use NAND2X1  NAND2X1_33
timestamp 1537603335
transform -1 0 876 0 1 305
box 0 0 24 100
use NOR2X1  NOR2X1_45
timestamp 1537603335
transform -1 0 900 0 1 305
box 0 0 24 100
use NOR2X1  NOR2X1_26
timestamp 1537603335
transform -1 0 924 0 1 305
box 0 0 24 100
use INVX1  INVX1_14
timestamp 1537603335
transform -1 0 940 0 1 305
box 0 0 16 100
use BUFX4  BUFX4_7
timestamp 1537603335
transform -1 0 972 0 1 305
box 0 0 32 100
use FILL  FILL_3_1_0
timestamp 1537603335
transform -1 0 980 0 1 305
box 0 0 8 100
use FILL  FILL_3_1_1
timestamp 1537603335
transform -1 0 988 0 1 305
box 0 0 8 100
use BUFX4  BUFX4_10
timestamp 1537603335
transform -1 0 1020 0 1 305
box 0 0 32 100
use OAI21X1  OAI21X1_7
timestamp 1537603335
transform 1 0 1020 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_4
timestamp 1537603335
transform 1 0 1052 0 1 305
box 0 0 32 100
use OAI21X1  OAI21X1_10
timestamp 1537603335
transform 1 0 1084 0 1 305
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_21
timestamp 1537603335
transform 1 0 1116 0 1 305
box 0 0 96 100
use AOI21X1  AOI21X1_13
timestamp 1537603335
transform 1 0 1212 0 1 305
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_7
timestamp 1537603335
transform 1 0 1244 0 1 305
box 0 0 96 100
use AOI21X1  AOI21X1_10
timestamp 1537603335
transform 1 0 1340 0 1 305
box 0 0 32 100
use NOR2X1  NOR2X1_20
timestamp 1537603335
transform -1 0 1396 0 1 305
box 0 0 24 100
use INVX1  INVX1_16
timestamp 1537603335
transform -1 0 1412 0 1 305
box 0 0 16 100
use BUFX2  BUFX2_20
timestamp 1537603335
transform 1 0 1412 0 1 305
box 0 0 24 100
use BUFX2  BUFX2_41
timestamp 1537603335
transform 1 0 1436 0 1 305
box 0 0 24 100
use FILL  FILL_4_1
timestamp 1537603335
transform 1 0 1460 0 1 305
box 0 0 8 100
use FILL  FILL_4_2
timestamp 1537603335
transform 1 0 1468 0 1 305
box 0 0 8 100
use FILL  FILL_4_3
timestamp 1537603335
transform 1 0 1476 0 1 305
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_44
timestamp 1537603335
transform -1 0 100 0 -1 305
box 0 0 96 100
use OAI21X1  OAI21X1_57
timestamp 1537603335
transform -1 0 132 0 -1 305
box 0 0 32 100
use NAND2X1  NAND2X1_43
timestamp 1537603335
transform -1 0 156 0 -1 305
box 0 0 24 100
use NOR3X1  NOR3X1_10
timestamp 1537603335
transform -1 0 220 0 -1 305
box 0 0 64 100
use OAI21X1  OAI21X1_47
timestamp 1537603335
transform 1 0 220 0 -1 305
box 0 0 32 100
use NOR2X1  NOR2X1_48
timestamp 1537603335
transform -1 0 276 0 -1 305
box 0 0 24 100
use NOR3X1  NOR3X1_20
timestamp 1537603335
transform -1 0 340 0 -1 305
box 0 0 64 100
use NOR2X1  NOR2X1_58
timestamp 1537603335
transform -1 0 364 0 -1 305
box 0 0 24 100
use AOI21X1  AOI21X1_25
timestamp 1537603335
transform 1 0 364 0 -1 305
box 0 0 32 100
use OAI22X1  OAI22X1_2
timestamp 1537603335
transform 1 0 396 0 -1 305
box 0 0 40 100
use NOR2X1  NOR2X1_57
timestamp 1537603335
transform -1 0 460 0 -1 305
box 0 0 24 100
use FILL  FILL_2_0_0
timestamp 1537603335
transform -1 0 468 0 -1 305
box 0 0 8 100
use FILL  FILL_2_0_1
timestamp 1537603335
transform -1 0 476 0 -1 305
box 0 0 8 100
use OAI22X1  OAI22X1_4
timestamp 1537603335
transform -1 0 516 0 -1 305
box 0 0 40 100
use NOR2X1  NOR2X1_60
timestamp 1537603335
transform -1 0 540 0 -1 305
box 0 0 24 100
use NAND3X1  NAND3X1_21
timestamp 1537603335
transform -1 0 572 0 -1 305
box 0 0 32 100
use OAI21X1  OAI21X1_51
timestamp 1537603335
transform -1 0 604 0 -1 305
box 0 0 32 100
use NOR2X1  NOR2X1_55
timestamp 1537603335
transform -1 0 628 0 -1 305
box 0 0 24 100
use NAND3X1  NAND3X1_25
timestamp 1537603335
transform -1 0 660 0 -1 305
box 0 0 32 100
use NOR3X1  NOR3X1_18
timestamp 1537603335
transform 1 0 660 0 -1 305
box 0 0 64 100
use INVX2  INVX2_10
timestamp 1537603335
transform 1 0 724 0 -1 305
box 0 0 16 100
use OAI21X1  OAI21X1_46
timestamp 1537603335
transform -1 0 772 0 -1 305
box 0 0 32 100
use NOR2X1  NOR2X1_42
timestamp 1537603335
transform -1 0 796 0 -1 305
box 0 0 24 100
use AND2X2  AND2X2_15
timestamp 1537603335
transform 1 0 796 0 -1 305
box 0 0 32 100
use INVX1  INVX1_35
timestamp 1537603335
transform -1 0 844 0 -1 305
box 0 0 16 100
use NAND2X1  NAND2X1_39
timestamp 1537603335
transform -1 0 868 0 -1 305
box 0 0 24 100
use INVX2  INVX2_5
timestamp 1537603335
transform 1 0 868 0 -1 305
box 0 0 16 100
use DFFPOSX1  DFFPOSX1_11
timestamp 1537603335
transform 1 0 884 0 -1 305
box 0 0 96 100
use FILL  FILL_2_1_0
timestamp 1537603335
transform 1 0 980 0 -1 305
box 0 0 8 100
use FILL  FILL_2_1_1
timestamp 1537603335
transform 1 0 988 0 -1 305
box 0 0 8 100
use BUFX2  BUFX2_26
timestamp 1537603335
transform 1 0 996 0 -1 305
box 0 0 24 100
use BUFX2  BUFX2_52
timestamp 1537603335
transform 1 0 1020 0 -1 305
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_17
timestamp 1537603335
transform -1 0 1140 0 -1 305
box 0 0 96 100
use INVX1  INVX1_20
timestamp 1537603335
transform 1 0 1140 0 -1 305
box 0 0 16 100
use NOR2X1  NOR2X1_32
timestamp 1537603335
transform 1 0 1156 0 -1 305
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_8
timestamp 1537603335
transform 1 0 1180 0 -1 305
box 0 0 96 100
use NOR2X1  NOR2X1_23
timestamp 1537603335
transform -1 0 1300 0 -1 305
box 0 0 24 100
use AOI21X1  AOI21X1_12
timestamp 1537603335
transform 1 0 1300 0 -1 305
box 0 0 32 100
use NOR2X1  NOR2X1_22
timestamp 1537603335
transform -1 0 1356 0 -1 305
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_5
timestamp 1537603335
transform 1 0 1356 0 -1 305
box 0 0 96 100
use BUFX2  BUFX2_23
timestamp 1537603335
transform 1 0 1452 0 -1 305
box 0 0 24 100
use FILL  FILL_3_1
timestamp 1537603335
transform -1 0 1484 0 -1 305
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_1
timestamp 1537603335
transform -1 0 100 0 1 105
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_46
timestamp 1537603335
transform -1 0 196 0 1 105
box 0 0 96 100
use NAND3X1  NAND3X1_24
timestamp 1537603335
transform -1 0 228 0 1 105
box 0 0 32 100
use INVX1  INVX1_31
timestamp 1537603335
transform -1 0 244 0 1 105
box 0 0 16 100
use NAND3X1  NAND3X1_16
timestamp 1537603335
transform 1 0 244 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_47
timestamp 1537603335
transform 1 0 276 0 1 105
box 0 0 24 100
use NAND2X1  NAND2X1_42
timestamp 1537603335
transform 1 0 300 0 1 105
box 0 0 24 100
use OAI21X1  OAI21X1_56
timestamp 1537603335
transform -1 0 356 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_44
timestamp 1537603335
transform 1 0 356 0 1 105
box 0 0 24 100
use INVX1  INVX1_30
timestamp 1537603335
transform -1 0 396 0 1 105
box 0 0 16 100
use NAND2X1  NAND2X1_31
timestamp 1537603335
transform -1 0 420 0 1 105
box 0 0 24 100
use NAND3X1  NAND3X1_22
timestamp 1537603335
transform 1 0 420 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_43
timestamp 1537603335
transform -1 0 476 0 1 105
box 0 0 24 100
use FILL  FILL_1_0_0
timestamp 1537603335
transform 1 0 476 0 1 105
box 0 0 8 100
use FILL  FILL_1_0_1
timestamp 1537603335
transform 1 0 484 0 1 105
box 0 0 8 100
use OAI22X1  OAI22X1_3
timestamp 1537603335
transform 1 0 492 0 1 105
box 0 0 40 100
use OAI21X1  OAI21X1_48
timestamp 1537603335
transform -1 0 564 0 1 105
box 0 0 32 100
use INVX2  INVX2_13
timestamp 1537603335
transform 1 0 564 0 1 105
box 0 0 16 100
use AOI21X1  AOI21X1_23
timestamp 1537603335
transform 1 0 580 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_52
timestamp 1537603335
transform -1 0 636 0 1 105
box 0 0 24 100
use NAND2X1  NAND2X1_44
timestamp 1537603335
transform 1 0 636 0 1 105
box 0 0 24 100
use NOR2X1  NOR2X1_54
timestamp 1537603335
transform -1 0 684 0 1 105
box 0 0 24 100
use INVX1  INVX1_33
timestamp 1537603335
transform 1 0 684 0 1 105
box 0 0 16 100
use NAND2X1  NAND2X1_40
timestamp 1537603335
transform -1 0 724 0 1 105
box 0 0 24 100
use NOR3X1  NOR3X1_19
timestamp 1537603335
transform 1 0 724 0 1 105
box 0 0 64 100
use NOR3X1  NOR3X1_15
timestamp 1537603335
transform 1 0 788 0 1 105
box 0 0 64 100
use NOR3X1  NOR3X1_17
timestamp 1537603335
transform 1 0 852 0 1 105
box 0 0 64 100
use NOR2X1  NOR2X1_5
timestamp 1537603335
transform -1 0 940 0 1 105
box 0 0 24 100
use NOR2X1  NOR2X1_6
timestamp 1537603335
transform -1 0 964 0 1 105
box 0 0 24 100
use NAND2X1  NAND2X1_4
timestamp 1537603335
transform -1 0 988 0 1 105
box 0 0 24 100
use FILL  FILL_1_1_0
timestamp 1537603335
transform 1 0 988 0 1 105
box 0 0 8 100
use FILL  FILL_1_1_1
timestamp 1537603335
transform 1 0 996 0 1 105
box 0 0 8 100
use AOI21X1  AOI21X1_7
timestamp 1537603335
transform 1 0 1004 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_17
timestamp 1537603335
transform 1 0 1036 0 1 105
box 0 0 24 100
use NOR2X1  NOR2X1_24
timestamp 1537603335
transform 1 0 1060 0 1 105
box 0 0 24 100
use AOI21X1  AOI21X1_14
timestamp 1537603335
transform -1 0 1116 0 1 105
box 0 0 32 100
use BUFX4  BUFX4_16
timestamp 1537603335
transform -1 0 1148 0 1 105
box 0 0 32 100
use BUFX4  BUFX4_13
timestamp 1537603335
transform 1 0 1148 0 1 105
box 0 0 32 100
use BUFX4  BUFX4_22
timestamp 1537603335
transform -1 0 1212 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_30
timestamp 1537603335
transform -1 0 1236 0 1 105
box 0 0 24 100
use INVX1  INVX1_18
timestamp 1537603335
transform -1 0 1252 0 1 105
box 0 0 16 100
use DFFPOSX1  DFFPOSX1_15
timestamp 1537603335
transform -1 0 1348 0 1 105
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_27
timestamp 1537603335
transform 1 0 1348 0 1 105
box 0 0 96 100
use BUFX4  BUFX4_21
timestamp 1537603335
transform 1 0 1444 0 1 105
box 0 0 32 100
use FILL  FILL_2_1
timestamp 1537603335
transform 1 0 1476 0 1 105
box 0 0 8 100
use BUFX2  BUFX2_60
timestamp 1537603335
transform -1 0 28 0 -1 105
box 0 0 24 100
use INVX2  INVX2_12
timestamp 1537603335
transform 1 0 28 0 -1 105
box 0 0 16 100
use AOI21X1  AOI21X1_24
timestamp 1537603335
transform 1 0 44 0 -1 105
box 0 0 32 100
use NOR2X1  NOR2X1_56
timestamp 1537603335
transform 1 0 76 0 -1 105
box 0 0 24 100
use NAND2X1  NAND2X1_35
timestamp 1537603335
transform -1 0 124 0 -1 105
box 0 0 24 100
use NOR3X1  NOR3X1_9
timestamp 1537603335
transform -1 0 188 0 -1 105
box 0 0 64 100
use NOR2X1  NOR2X1_46
timestamp 1537603335
transform -1 0 212 0 -1 105
box 0 0 24 100
use NOR3X1  NOR3X1_13
timestamp 1537603335
transform 1 0 212 0 -1 105
box 0 0 64 100
use INVX2  INVX2_11
timestamp 1537603335
transform 1 0 276 0 -1 105
box 0 0 16 100
use OAI21X1  OAI21X1_53
timestamp 1537603335
transform 1 0 292 0 -1 105
box 0 0 32 100
use OAI21X1  OAI21X1_52
timestamp 1537603335
transform -1 0 356 0 -1 105
box 0 0 32 100
use NOR3X1  NOR3X1_11
timestamp 1537603335
transform 1 0 356 0 -1 105
box 0 0 64 100
use NAND3X1  NAND3X1_15
timestamp 1537603335
transform 1 0 420 0 -1 105
box 0 0 32 100
use NOR2X1  NOR2X1_53
timestamp 1537603335
transform -1 0 476 0 -1 105
box 0 0 24 100
use FILL  FILL_0_0_0
timestamp 1537603335
transform 1 0 476 0 -1 105
box 0 0 8 100
use FILL  FILL_0_0_1
timestamp 1537603335
transform 1 0 484 0 -1 105
box 0 0 8 100
use OAI21X1  OAI21X1_54
timestamp 1537603335
transform 1 0 492 0 -1 105
box 0 0 32 100
use NOR3X1  NOR3X1_16
timestamp 1537603335
transform 1 0 524 0 -1 105
box 0 0 64 100
use OAI21X1  OAI21X1_55
timestamp 1537603335
transform 1 0 588 0 -1 105
box 0 0 32 100
use NAND2X1  NAND2X1_41
timestamp 1537603335
transform -1 0 644 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_34
timestamp 1537603335
transform 1 0 644 0 -1 105
box 0 0 24 100
use NAND3X1  NAND3X1_23
timestamp 1537603335
transform 1 0 668 0 -1 105
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_45
timestamp 1537603335
transform -1 0 796 0 -1 105
box 0 0 96 100
use BUFX2  BUFX2_50
timestamp 1537603335
transform -1 0 820 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_51
timestamp 1537603335
transform -1 0 844 0 -1 105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_2
timestamp 1537603335
transform 1 0 844 0 -1 105
box 0 0 96 100
use BUFX2  BUFX2_17
timestamp 1537603335
transform 1 0 940 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_24
timestamp 1537603335
transform 1 0 964 0 -1 105
box 0 0 24 100
use FILL  FILL_0_1_0
timestamp 1537603335
transform -1 0 996 0 -1 105
box 0 0 8 100
use FILL  FILL_0_1_1
timestamp 1537603335
transform -1 0 1004 0 -1 105
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_9
timestamp 1537603335
transform -1 0 1100 0 -1 105
box 0 0 96 100
use BUFX2  BUFX2_32
timestamp 1537603335
transform 1 0 1100 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_38
timestamp 1537603335
transform 1 0 1124 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_66
timestamp 1537603335
transform 1 0 1148 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_72
timestamp 1537603335
transform 1 0 1172 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_46
timestamp 1537603335
transform 1 0 1196 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_67
timestamp 1537603335
transform 1 0 1220 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_30
timestamp 1537603335
transform 1 0 1244 0 -1 105
box 0 0 24 100
use XOR2X1  XOR2X1_1
timestamp 1537603335
transform 1 0 1268 0 -1 105
box 0 0 56 100
use BUFX2  BUFX2_33
timestamp 1537603335
transform 1 0 1324 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_68
timestamp 1537603335
transform -1 0 1372 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_40
timestamp 1537603335
transform 1 0 1372 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_43
timestamp 1537603335
transform 1 0 1396 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_42
timestamp 1537603335
transform 1 0 1420 0 -1 105
box 0 0 24 100
use NAND2X1  NAND2X1_16
timestamp 1537603335
transform 1 0 1444 0 -1 105
box 0 0 24 100
use FILL  FILL_1_1
timestamp 1537603335
transform -1 0 1476 0 -1 105
box 0 0 8 100
use FILL  FILL_1_2
timestamp 1537603335
transform -1 0 1484 0 -1 105
box 0 0 8 100
<< labels >>
rlabel metal6 s 472 -30 488 -22 8 vdd
port 0 nsew
rlabel metal6 s 976 -30 992 -22 8 gnd
port 1 nsew
rlabel metal3 s -24 460 -24 460 4 clk
port 2 nsew
rlabel metal2 s 920 -20 920 -20 8 INPD<0>
port 3 nsew
rlabel metal2 s 1120 1230 1120 1230 6 INPD<1>
port 4 nsew
rlabel metal2 s 1184 1230 1184 1230 6 INPD<2>
port 5 nsew
rlabel metal3 s 1512 780 1512 780 6 INPD<3>
port 6 nsew
rlabel metal3 s 1512 760 1512 760 6 INPD<4>
port 7 nsew
rlabel metal3 s 1512 720 1512 720 6 INPD<5>
port 8 nsew
rlabel metal3 s 1512 960 1512 960 6 INPD<6>
port 9 nsew
rlabel metal3 s 1512 530 1512 530 6 INPD<7>
port 10 nsew
rlabel metal2 s 1080 -20 1080 -20 8 INPD<8>
port 11 nsew
rlabel metal2 s 984 1230 984 1230 6 INPD<9>
port 12 nsew
rlabel metal2 s 464 1230 464 1230 6 INPD<10>
port 13 nsew
rlabel metal2 s 1040 1230 1040 1230 6 INPD<11>
port 14 nsew
rlabel metal3 s -24 1180 -24 1180 4 INPD<12>
port 15 nsew
rlabel metal3 s -24 1130 -24 1130 4 INPD<13>
port 16 nsew
rlabel metal2 s 40 1230 40 1230 6 INPD<14>
port 17 nsew
rlabel metal3 s 1512 510 1512 510 6 INPD<15>
port 18 nsew
rlabel metal2 s 888 -20 888 -20 8 RDATA<0>
port 19 nsew
rlabel metal2 s 1096 1230 1096 1230 6 RDATA<1>
port 20 nsew
rlabel metal3 s 1512 740 1512 740 6 RDATA<2>
port 21 nsew
rlabel metal3 s 1512 600 1512 600 6 RDATA<3>
port 22 nsew
rlabel metal3 s 1512 660 1512 660 6 RDATA<4>
port 23 nsew
rlabel metal3 s 1512 160 1512 160 6 RDATA<5>
port 24 nsew
rlabel metal2 s 1136 1230 1136 1230 6 RDATA<6>
port 25 nsew
rlabel metal3 s 1512 680 1512 680 6 RDATA<7>
port 26 nsew
rlabel metal2 s 424 -20 424 -20 8 RF
port 27 nsew
rlabel metal3 s -24 80 -24 80 4 WF
port 28 nsew
rlabel metal2 s 368 -20 368 -20 8 NEXTOP<0>
port 29 nsew
rlabel metal2 s 720 -20 720 -20 8 NEXTOP<1>
port 30 nsew
rlabel metal2 s 616 -20 616 -20 8 NEXTOP<2>
port 31 nsew
rlabel metal2 s 1056 1230 1056 1230 6 IR
port 32 nsew
rlabel metal2 s 1344 -20 1344 -20 8 OW
port 33 nsew
rlabel metal2 s 960 -20 960 -20 8 OUTPD<0>
port 34 nsew
rlabel metal2 s 1232 1230 1232 1230 6 OUTPD<1>
port 35 nsew
rlabel metal2 s 1256 1230 1256 1230 6 OUTPD<2>
port 36 nsew
rlabel metal3 s 1512 380 1512 380 6 OUTPD<3>
port 37 nsew
rlabel metal3 s 1512 460 1512 460 6 OUTPD<4>
port 38 nsew
rlabel metal3 s 1512 580 1512 580 6 OUTPD<5>
port 39 nsew
rlabel metal3 s 1512 260 1512 260 6 OUTPD<6>
port 40 nsew
rlabel metal2 s 984 -20 984 -20 8 OUTPD<7>
port 41 nsew
rlabel metal3 s -24 360 -24 360 4 OUTPD<8>
port 42 nsew
rlabel metal2 s 1024 -20 1024 -20 8 OUTPD<9>
port 43 nsew
rlabel metal3 s -24 1060 -24 1060 4 OUTPD<10>
port 44 nsew
rlabel metal2 s 1376 1230 1376 1230 6 OUTPD<11>
port 45 nsew
rlabel metal3 s -24 580 -24 580 4 OUTPD<12>
port 46 nsew
rlabel metal2 s 1264 -20 1264 -20 8 OUTPD<13>
port 47 nsew
rlabel metal2 s 872 1230 872 1230 6 OUTPD<14>
port 48 nsew
rlabel metal2 s 1120 -20 1120 -20 8 OUTPD<15>
port 49 nsew
rlabel metal3 s -24 60 -24 60 4 reset
port 50 nsew
rlabel metal2 s 800 -20 800 -20 8 RD
port 51 nsew
rlabel metal2 s 824 -20 824 -20 8 WD
port 52 nsew
rlabel metal2 s 1040 -20 1040 -20 8 WDATA<0>
port 53 nsew
rlabel metal2 s 952 1230 952 1230 6 WDATA<1>
port 54 nsew
rlabel metal2 s 1000 1230 1000 1230 6 WDATA<2>
port 55 nsew
rlabel metal3 s 1512 560 1512 560 6 WDATA<3>
port 56 nsew
rlabel metal3 s 1512 800 1512 800 6 WDATA<4>
port 57 nsew
rlabel metal2 s 1080 1230 1080 1230 6 WDATA<5>
port 58 nsew
rlabel metal3 s 1512 980 1512 980 6 WDATA<6>
port 59 nsew
rlabel metal3 s 1512 860 1512 860 6 WDATA<7>
port 60 nsew
rlabel metal3 s -24 760 -24 760 4 DP<0>
port 61 nsew
rlabel metal3 s -24 980 -24 980 4 DP<1>
port 62 nsew
rlabel metal3 s -24 960 -24 960 4 DP<2>
port 63 nsew
rlabel metal3 s -24 660 -24 660 4 DP<3>
port 64 nsew
rlabel metal2 s 632 -20 632 -20 8 DP<4>
port 65 nsew
rlabel metal2 s 592 -20 592 -20 8 DP<5>
port 66 nsew
rlabel metal2 s 848 1230 848 1230 6 DP<6>
port 67 nsew
rlabel metal2 s 616 1230 616 1230 6 DP<7>
port 68 nsew
rlabel metal3 s -24 860 -24 860 4 DP<8>
port 69 nsew
rlabel metal2 s 480 1230 480 1230 6 DP<9>
port 70 nsew
rlabel metal2 s 168 1230 168 1230 6 DP<10>
port 71 nsew
rlabel metal2 s 104 1230 104 1230 6 DP<11>
port 72 nsew
rlabel metal2 s 824 1230 824 1230 6 DP<12>
port 73 nsew
rlabel metal2 s 704 1230 704 1230 6 DP<13>
port 74 nsew
rlabel metal2 s 216 1230 216 1230 6 DP<14>
port 75 nsew
rlabel metal2 s 664 -20 664 -20 8 PCDELTA<0>
port 76 nsew
rlabel metal3 s -24 560 -24 560 4 PCDELTA<1>
port 77 nsew
rlabel metal2 s 1448 1230 1448 1230 6 PCDELTA<2>
port 78 nsew
rlabel metal2 s 912 1230 912 1230 6 PCDELTA<3>
port 79 nsew
rlabel metal2 s 1144 -20 1144 -20 8 PCDELTA<4>
port 80 nsew
rlabel metal2 s 936 1230 936 1230 6 PCDELTA<5>
port 81 nsew
rlabel metal2 s 1392 -20 1392 -20 8 PCDELTA<6>
port 82 nsew
rlabel metal3 s 1512 360 1512 360 6 PCDELTA<7>
port 83 nsew
rlabel metal2 s 1440 -20 1440 -20 8 PCDELTA<8>
port 84 nsew
rlabel metal2 s 1416 -20 1416 -20 8 PCDELTA<9>
port 85 nsew
rlabel metal3 s 1512 1000 1512 1000 6 PCDELTA<10>
port 86 nsew
rlabel metal2 s 1424 1230 1424 1230 6 PCDELTA<11>
port 87 nsew
rlabel metal2 s 1216 -20 1216 -20 8 PCDELTA<12>
port 88 nsew
rlabel metal3 s 1512 700 1512 700 6 PCDELTA<13>
port 89 nsew
rlabel metal3 s 1512 1160 1512 1160 6 PCDELTA<14>
port 90 nsew
rlabel metal2 s 896 1230 896 1230 6 PCDELTA<15>
port 91 nsew
<< end >>
