* XSpice netlist created from SPICE and liberty sources by spi2xspice.py
*SPICE netlist created from BLIF module BFCPU by blif2BSpice
.subckt BFCPU a_vdd a_gnd a_clk a_INPD_0_ a_INPD_1_ a_INPD_2_ a_INPD_3_ a_INPD_4_ a_INPD_5_ a_INPD_6_ a_INPD_7_ a_INPD_8_ a_INPD_9_ a_INPD_10_ a_INPD_11_ a_INPD_12_ a_INPD_13_ a_INPD_14_ a_INPD_15_ a_RDATA_0_ a_RDATA_1_ a_RDATA_2_ a_RDATA_3_ a_RDATA_4_ a_RDATA_5_ a_RDATA_6_ a_RDATA_7_ a_RF a_WF a_NEXTOP_0_ a_NEXTOP_1_ a_NEXTOP_2_ a_IR a_OW a_OUTPD_0_ a_OUTPD_1_ a_OUTPD_2_ a_OUTPD_3_ a_OUTPD_4_ a_OUTPD_5_ a_OUTPD_6_ a_OUTPD_7_ a_OUTPD_8_ a_OUTPD_9_ a_OUTPD_10_ a_OUTPD_11_ a_OUTPD_12_ a_OUTPD_13_ a_OUTPD_14_ a_OUTPD_15_ a_reset a_RD a_WD a_WDATA_0_ a_WDATA_1_ a_WDATA_2_ a_WDATA_3_ a_WDATA_4_ a_WDATA_5_ a_WDATA_6_ a_WDATA_7_ a_DP_0_ a_DP_1_ a_DP_2_ a_DP_3_ a_DP_4_ a_DP_5_ a_DP_6_ a_DP_7_ a_DP_8_ a_DP_9_ a_DP_10_ a_DP_11_ a_DP_12_ a_DP_13_ a_DP_14_ a_PCDELTA_0_ a_PCDELTA_1_ a_PCDELTA_2_ a_PCDELTA_3_ a_PCDELTA_4_ a_PCDELTA_5_ a_PCDELTA_6_ a_PCDELTA_7_ a_PCDELTA_8_ a_PCDELTA_9_ a_PCDELTA_10_ a_PCDELTA_11_ a_PCDELTA_12_ a_PCDELTA_13_ a_PCDELTA_14_ a_PCDELTA_15_
ABUFX4_1 [DC1.SGN] DC1.SGN_bF$buf5 d_lut_BUFX4
ABUFX4_2 [DC1.SGN] DC1.SGN_bF$buf4 d_lut_BUFX4
ABUFX4_3 [DC1.SGN] DC1.SGN_bF$buf3 d_lut_BUFX4
ABUFX4_4 [DC1.SGN] DC1.SGN_bF$buf2 d_lut_BUFX4
ABUFX4_5 [DC1.SGN] DC1.SGN_bF$buf1 d_lut_BUFX4
ABUFX4_6 [DC1.SGN] DC1.SGN_bF$buf0 d_lut_BUFX4
ABUFX4_7 [clk] clk_bF$buf5 d_lut_BUFX4
ABUFX4_8 [clk] clk_bF$buf4 d_lut_BUFX4
ABUFX4_9 [clk] clk_bF$buf3 d_lut_BUFX4
ABUFX4_10 [clk] clk_bF$buf2 d_lut_BUFX4
ABUFX4_11 [clk] clk_bF$buf1 d_lut_BUFX4
ABUFX4_12 [clk] clk_bF$buf0 d_lut_BUFX4
ABUFX4_13 [_119_] _119__bF$buf4 d_lut_BUFX4
ABUFX4_14 [_119_] _119__bF$buf3 d_lut_BUFX4
ABUFX4_15 [_119_] _119__bF$buf2 d_lut_BUFX4
ABUFX4_16 [_119_] _119__bF$buf1 d_lut_BUFX4
ABUFX4_17 [_119_] _119__bF$buf0 d_lut_BUFX4
ABUFX4_18 [OPC1.PCDELTA_15_] OPC1.PCDELTA_15_bF$buf4 d_lut_BUFX4
ABUFX4_19 [OPC1.PCDELTA_15_] OPC1.PCDELTA_15_bF$buf3 d_lut_BUFX4
ABUFX4_20 [OPC1.PCDELTA_15_] OPC1.PCDELTA_15_bF$buf2 d_lut_BUFX4
ABUFX4_21 [OPC1.PCDELTA_15_] OPC1.PCDELTA_15_bF$buf1 d_lut_BUFX4
ABUFX4_22 [OPC1.PCDELTA_15_] OPC1.PCDELTA_15_bF$buf0 d_lut_BUFX4
AINVX1_1 [OPC1.INST_3_] _0_ d_lut_INVX1
ANAND2X1_1 [OPC1.INST_2_ _0_] _1_ d_lut_NAND2X1
AOR2X2_1 [OPC1.INST_1_ DC1.SGN_bF$buf5] _2_ d_lut_OR2X2
ANOR2X1_1 [_2_ _1_] DC1.OUTP d_lut_NOR2X1
AINVX1_2 [OPC1.INST_2_] _3_ d_lut_INVX1
ANAND2X1_2 [OPC1.INST_1_ _3_] _4_ d_lut_NAND2X1
ANOR2X1_2 [OPC1.INST_3_ _4_] DC1.DOP d_lut_NOR2X1
ANOR2X1_3 [OPC1.INST_1_ OPC1.INST_3_] _5_ d_lut_NOR2X1
AAND2X2_1 [_5_ _3_] DPC1.DPOP d_lut_AND2X2
ANAND2X1_3 [DC1.SGN_bF$buf4 OPC1.INST_3_] _6_ d_lut_NAND2X1
ANOR2X1_4 [_6_ _4_] DC1.LD d_lut_NOR2X1
ANAND2X1_4 [OPC1.INST_3_ OPC1.INST_2_] _7_ d_lut_NAND2X1
ANOR2X1_5 [_7_ _2_] _10_ d_lut_NOR2X1
AINVX1_3 [OPC1.INST_1_] _8_ d_lut_INVX1
ANAND2X1_5 [DC1.SGN_bF$buf3 _8_] _9_ d_lut_NAND2X1
ANOR2X1_6 [_7_ _9_] _11_ d_lut_NOR2X1
ANOR2X1_7 [_1_ _9_] DC1.INP d_lut_NOR2X1
ABUFX2_1 [DPC1.DP_0_] DP_0_ d_lut_BUFX2
ABUFX2_2 [DPC1.DP_1_] DP_1_ d_lut_BUFX2
ABUFX2_3 [DPC1.DP_2_] DP_2_ d_lut_BUFX2
ABUFX2_4 [DPC1.DP_3_] DP_3_ d_lut_BUFX2
ABUFX2_5 [DPC1.DP_4_] DP_4_ d_lut_BUFX2
ABUFX2_6 [DPC1.DP_5_] DP_5_ d_lut_BUFX2
ABUFX2_7 [DPC1.DP_6_] DP_6_ d_lut_BUFX2
ABUFX2_8 [DPC1.DP_7_] DP_7_ d_lut_BUFX2
ABUFX2_9 [DPC1.DP_8_] DP_8_ d_lut_BUFX2
ABUFX2_10 [DPC1.DP_9_] DP_9_ d_lut_BUFX2
ABUFX2_11 [DPC1.DP_10_] DP_10_ d_lut_BUFX2
ABUFX2_12 [DPC1.DP_11_] DP_11_ d_lut_BUFX2
ABUFX2_13 [DPC1.DP_12_] DP_12_ d_lut_BUFX2
ABUFX2_14 [DPC1.DP_13_] DP_13_ d_lut_BUFX2
ABUFX2_15 [DPC1.DP_14_] DP_14_ d_lut_BUFX2
ABUFX2_16 [DC1.IR] IR d_lut_BUFX2
ABUFX2_17 [DC1.OUTPD_0_] OUTPD_0_ d_lut_BUFX2
ABUFX2_18 [DC1.OUTPD_1_] OUTPD_1_ d_lut_BUFX2
ABUFX2_19 [DC1.OUTPD_2_] OUTPD_2_ d_lut_BUFX2
ABUFX2_20 [DC1.OUTPD_3_] OUTPD_3_ d_lut_BUFX2
ABUFX2_21 [DC1.OUTPD_4_] OUTPD_4_ d_lut_BUFX2
ABUFX2_22 [DC1.OUTPD_5_] OUTPD_5_ d_lut_BUFX2
ABUFX2_23 [DC1.OUTPD_6_] OUTPD_6_ d_lut_BUFX2
ABUFX2_24 [DC1.OUTPD_7_] OUTPD_7_ d_lut_BUFX2
ABUFX2_25 [DC1.OUTPD_8_] OUTPD_8_ d_lut_BUFX2
ABUFX2_26 [DC1.OUTPD_9_] OUTPD_9_ d_lut_BUFX2
ABUFX2_27 [DC1.OUTPD_10_] OUTPD_10_ d_lut_BUFX2
ABUFX2_28 [DC1.OUTPD_11_] OUTPD_11_ d_lut_BUFX2
ABUFX2_29 [DC1.OUTPD_12_] OUTPD_12_ d_lut_BUFX2
ABUFX2_30 [DC1.OUTPD_13_] OUTPD_13_ d_lut_BUFX2
ABUFX2_31 [DC1.OUTPD_14_] OUTPD_14_ d_lut_BUFX2
ABUFX2_32 [DC1.OUTPD_15_] OUTPD_15_ d_lut_BUFX2
ABUFX2_33 [DC1.OW] OW d_lut_BUFX2
ABUFX2_34 [OPC1.PCDELTA_0_] PCDELTA_0_ d_lut_BUFX2
ABUFX2_35 [OPC1.PCDELTA_15_bF$buf4] PCDELTA_1_ d_lut_BUFX2
ABUFX2_36 [OPC1.PCDELTA_15_bF$buf3] PCDELTA_2_ d_lut_BUFX2
ABUFX2_37 [OPC1.PCDELTA_15_bF$buf2] PCDELTA_3_ d_lut_BUFX2
ABUFX2_38 [OPC1.PCDELTA_15_bF$buf1] PCDELTA_4_ d_lut_BUFX2
ABUFX2_39 [OPC1.PCDELTA_15_bF$buf0] PCDELTA_5_ d_lut_BUFX2
ABUFX2_40 [OPC1.PCDELTA_15_bF$buf4] PCDELTA_6_ d_lut_BUFX2
ABUFX2_41 [OPC1.PCDELTA_15_bF$buf3] PCDELTA_7_ d_lut_BUFX2
ABUFX2_42 [OPC1.PCDELTA_15_bF$buf2] PCDELTA_8_ d_lut_BUFX2
ABUFX2_43 [OPC1.PCDELTA_15_bF$buf1] PCDELTA_9_ d_lut_BUFX2
ABUFX2_44 [OPC1.PCDELTA_15_bF$buf0] PCDELTA_10_ d_lut_BUFX2
ABUFX2_45 [OPC1.PCDELTA_15_bF$buf4] PCDELTA_11_ d_lut_BUFX2
ABUFX2_46 [OPC1.PCDELTA_15_bF$buf3] PCDELTA_12_ d_lut_BUFX2
ABUFX2_47 [OPC1.PCDELTA_15_bF$buf2] PCDELTA_13_ d_lut_BUFX2
ABUFX2_48 [OPC1.PCDELTA_15_bF$buf1] PCDELTA_14_ d_lut_BUFX2
ABUFX2_49 [OPC1.PCDELTA_15_bF$buf0] PCDELTA_15_ d_lut_BUFX2
ABUFX2_50 [_10_] RD d_lut_BUFX2
ABUFX2_51 [_11_] WD d_lut_BUFX2
ABUFX2_52 [DC1.WDATA_0_] WDATA_0_ d_lut_BUFX2
ABUFX2_53 [DC1.WDATA_1_] WDATA_1_ d_lut_BUFX2
ABUFX2_54 [DC1.WDATA_2_] WDATA_2_ d_lut_BUFX2
ABUFX2_55 [DC1.WDATA_3_] WDATA_3_ d_lut_BUFX2
ABUFX2_56 [DC1.WDATA_4_] WDATA_4_ d_lut_BUFX2
ABUFX2_57 [DC1.WDATA_5_] WDATA_5_ d_lut_BUFX2
ABUFX2_58 [DC1.WDATA_6_] WDATA_6_ d_lut_BUFX2
ABUFX2_59 [DC1.WDATA_7_] WDATA_7_ d_lut_BUFX2
ABUFX2_60 [_12_] reset d_lut_BUFX2
ADFFPOSX1_1 vdd clk_bF$buf5 NULL NULL _12_ NULL ddflop
AINVX4_1 [DC1.WDATA_2_] _107_ d_lut_INVX4
AINVX2_1 [DC1.WDATA_5_] _108_ d_lut_INVX2
ANOR2X1_8 [DC1.WDATA_3_ DC1.WDATA_4_] _109_ d_lut_NOR2X1
ANAND3X1_1 [_107_ _108_ _109_] _110_ d_lut_NAND3X1
AINVX2_2 [DC1.WDATA_7_] _111_ d_lut_INVX2
AINVX4_2 [DC1.WDATA_6_] _112_ d_lut_INVX4
ANOR2X1_9 [DC1.WDATA_1_ DC1.WDATA_0_] _113_ d_lut_NOR2X1
ANAND3X1_2 [_111_ _112_ _113_] _114_ d_lut_NAND3X1
ANOR2X1_10 [_110_ _114_] DC1.IZ d_lut_NOR2X1
AINVX2_3 [DC1.LD] _115_ d_lut_INVX2
ANAND2X1_6 [DC1.OUTP _115_] _116_ d_lut_NAND2X1
ANOR2X1_11 [DC1.INP DC1.DOP] _117_ d_lut_NOR2X1
AINVX1_4 [_117_] _118_ d_lut_INVX1
ANOR2X1_12 [_116_ _118_] _119_ d_lut_NOR2X1
AXOR2X1_1 [_119__bF$buf4 DC1.OW] _15_ d_lut_XOR2X1
AINVX2_4 [DC1.INP] _120_ d_lut_INVX2
ANOR2X1_13 [DC1.DOP _120_] _121_ d_lut_NOR2X1
AXOR2X1_2 [_121_ DC1.IR] _13_ d_lut_XOR2X1
AINVX2_5 [DC1.WDATA_0_] _122_ d_lut_INVX2
ANAND2X1_7 [_122_ _115_] _123_ d_lut_NAND2X1
AOAI21X1_1 [_115_ RDATA_0_ _123_] _124_ d_lut_OAI21X1
AAOI22X1_1 [_122_ DC1.DOP _121_ INPD_0_] _125_ d_lut_AOI22X1
AOAI21X1_2 [_118_ _124_ _125_] _16__0_ d_lut_OAI21X1
AAND2X2_2 [DC1.WDATA_1_ DC1.WDATA_0_] _126_ d_lut_AND2X2
ANOR2X1_14 [_113_ _126_] _127_ d_lut_NOR2X1
AXNOR2X1_1 [_127_ DC1.SGN_bF$buf2] _17_ d_lut_XNOR2X1
AINVX1_5 [DC1.WDATA_1_] _18_ d_lut_INVX1
ANAND2X1_8 [DC1.LD RDATA_1_] _19_ d_lut_NAND2X1
AOAI21X1_3 [_18_ DC1.LD _19_] _20_ d_lut_OAI21X1
AMUX2X1_1 [_20_ INPD_1_ _120_] _21_ d_lut_MUX2X1
AMUX2X1_2 [_17_ _21_ DC1.DOP] _16__1_ d_lut_MUX2X1
ANAND2X1_9 [DC1.LD RDATA_2_] _22_ d_lut_NAND2X1
AOAI21X1_4 [_107_ DC1.LD _22_] _23_ d_lut_OAI21X1
AMUX2X1_3 [_23_ INPD_2_ _120_] _24_ d_lut_MUX2X1
AMUX2X1_4 [_113_ _126_ DC1.SGN_bF$buf1] _25_ d_lut_MUX2X1
AAND2X2_3 [_25_ _107_] _26_ d_lut_AND2X2
AOAI21X1_5 [_25_ _107_ DC1.DOP] _27_ d_lut_OAI21X1
AOAI22X1_1 [DC1.DOP _24_ _26_ _27_] _16__2_ d_lut_OAI22X1
ANOR3X1_1 [DC1.WDATA_1_ DC1.WDATA_0_ DC1.WDATA_2_] _28_ d_lut_NOR3X1
ANAND2X1_10 [DC1.SGN_bF$buf0 _28_] _29_ d_lut_NAND2X1
ANAND2X1_11 [DC1.WDATA_2_ _126_] _30_ d_lut_NAND2X1
AOAI21X1_6 [_30_ DC1.SGN_bF$buf5 _29_] _31_ d_lut_OAI21X1
AAND2X2_4 [_31_ DC1.WDATA_3_] _32_ d_lut_AND2X2
AOAI21X1_7 [_31_ DC1.WDATA_3_ DC1.DOP] _33_ d_lut_OAI21X1
AINVX1_6 [DC1.WDATA_3_] _34_ d_lut_INVX1
ANAND2X1_12 [DC1.LD RDATA_3_] _35_ d_lut_NAND2X1
AOAI21X1_8 [_34_ DC1.LD _35_] _36_ d_lut_OAI21X1
AINVX1_7 [INPD_3_] _37_ d_lut_INVX1
AAOI21X1_1 [DC1.INP _37_ DC1.DOP] _38_ d_lut_AOI21X1
AOAI21X1_9 [_36_ DC1.INP _38_] _39_ d_lut_OAI21X1
AOAI21X1_10 [_32_ _33_ _39_] _16__3_ d_lut_OAI21X1
AINVX2_6 [DC1.WDATA_4_] _40_ d_lut_INVX2
AINVX1_8 [DC1.SGN_bF$buf4] _41_ d_lut_INVX1
ANAND2X1_13 [DC1.WDATA_1_ DC1.WDATA_0_] _42_ d_lut_NAND2X1
ANAND2X1_14 [DC1.WDATA_3_ DC1.WDATA_2_] _43_ d_lut_NAND2X1
ANOR2X1_15 [_42_ _43_] _44_ d_lut_NOR2X1
ANOR2X1_16 [DC1.WDATA_3_ _41_] _45_ d_lut_NOR2X1
AAOI22X1_2 [_28_ _45_ _44_ _41_] _46_ d_lut_AOI22X1
AAND2X2_5 [_46_ _40_] _47_ d_lut_AND2X2
AOAI21X1_11 [_46_ _40_ DC1.DOP] _48_ d_lut_OAI21X1
ANAND2X1_15 [DC1.LD RDATA_4_] _49_ d_lut_NAND2X1
AOAI21X1_12 [_40_ DC1.LD _49_] _50_ d_lut_OAI21X1
AINVX1_9 [INPD_4_] _51_ d_lut_INVX1
AAOI21X1_2 [DC1.INP _51_ DC1.DOP] _52_ d_lut_AOI21X1
AOAI21X1_13 [_50_ DC1.INP _52_] _53_ d_lut_OAI21X1
AOAI21X1_14 [_47_ _48_ _53_] _16__4_ d_lut_OAI21X1
ANAND3X1_3 [DC1.SGN_bF$buf3 _109_ _28_] _54_ d_lut_NAND3X1
AAND2X2_6 [DC1.WDATA_3_ DC1.WDATA_2_] _55_ d_lut_AND2X2
ANAND3X1_4 [DC1.WDATA_4_ _126_ _55_] _56_ d_lut_NAND3X1
AOAI21X1_15 [_56_ DC1.SGN_bF$buf2 _54_] _57_ d_lut_OAI21X1
AAND2X2_7 [_57_ DC1.WDATA_5_] _58_ d_lut_AND2X2
AOAI21X1_16 [_57_ DC1.WDATA_5_ DC1.DOP] _59_ d_lut_OAI21X1
ANAND2X1_16 [DC1.LD RDATA_5_] _60_ d_lut_NAND2X1
AOAI21X1_17 [_108_ DC1.LD _60_] _61_ d_lut_OAI21X1
AINVX1_10 [INPD_5_] _62_ d_lut_INVX1
AAOI21X1_3 [DC1.INP _62_ DC1.DOP] _63_ d_lut_AOI21X1
AOAI21X1_18 [_61_ DC1.INP _63_] _64_ d_lut_OAI21X1
AOAI21X1_19 [_58_ _59_ _64_] _16__5_ d_lut_OAI21X1
ANOR3X1_2 [DC1.WDATA_3_ DC1.WDATA_5_ DC1.WDATA_4_] _65_ d_lut_NOR3X1
ANAND3X1_5 [DC1.SGN_bF$buf1 _28_ _65_] _66_ d_lut_NAND3X1
AAND2X2_8 [DC1.WDATA_5_ DC1.WDATA_4_] _67_ d_lut_AND2X2
ANAND3X1_6 [_126_ _55_ _67_] _68_ d_lut_NAND3X1
AOAI21X1_20 [_68_ DC1.SGN_bF$buf0 _66_] _69_ d_lut_OAI21X1
AAND2X2_9 [_69_ DC1.WDATA_6_] _70_ d_lut_AND2X2
AOAI21X1_21 [_69_ DC1.WDATA_6_ DC1.DOP] _71_ d_lut_OAI21X1
ANAND2X1_17 [DC1.LD RDATA_6_] _72_ d_lut_NAND2X1
AOAI21X1_22 [_112_ DC1.LD _72_] _73_ d_lut_OAI21X1
AINVX1_11 [INPD_6_] _74_ d_lut_INVX1
AAOI21X1_4 [DC1.INP _74_ DC1.DOP] _75_ d_lut_AOI21X1
AOAI21X1_23 [_73_ DC1.INP _75_] _76_ d_lut_OAI21X1
AOAI21X1_24 [_70_ _71_ _76_] _16__6_ d_lut_OAI21X1
ANAND2X1_18 [DC1.WDATA_5_ DC1.WDATA_4_] _77_ d_lut_NAND2X1
ANOR3X1_3 [_42_ _43_ _77_] _78_ d_lut_NOR3X1
ANAND3X1_7 [DC1.WDATA_7_ DC1.WDATA_6_ _78_] _79_ d_lut_NAND3X1
AOAI21X1_25 [_68_ _112_ _111_] _80_ d_lut_OAI21X1
AAOI21X1_5 [_79_ _80_ DC1.SGN_bF$buf5] _81_ d_lut_AOI21X1
ANAND3X1_8 [_112_ _28_ _65_] _82_ d_lut_NAND3X1
AAND2X2_10 [_82_ DC1.WDATA_7_] _83_ d_lut_AND2X2
AOAI21X1_26 [_110_ _114_ DC1.SGN_bF$buf4] _84_ d_lut_OAI21X1
AOAI21X1_27 [_83_ _84_ DC1.DOP] _85_ d_lut_OAI21X1
ANAND2X1_19 [DC1.LD RDATA_7_] _86_ d_lut_NAND2X1
AOAI21X1_28 [_111_ DC1.LD _86_] _87_ d_lut_OAI21X1
AINVX1_12 [INPD_7_] _88_ d_lut_INVX1
AAOI21X1_6 [DC1.INP _88_ DC1.DOP] _89_ d_lut_AOI21X1
AOAI21X1_29 [_87_ DC1.INP _89_] _90_ d_lut_OAI21X1
AOAI21X1_30 [_85_ _81_ _90_] _16__7_ d_lut_OAI21X1
ANOR2X1_17 [DC1.OUTPD_0_ _119__bF$buf3] _91_ d_lut_NOR2X1
AAOI21X1_7 [_122_ _119__bF$buf2 _91_] _14__0_ d_lut_AOI21X1
ANOR2X1_18 [DC1.OUTPD_1_ _119__bF$buf1] _92_ d_lut_NOR2X1
AAOI21X1_8 [_18_ _119__bF$buf0 _92_] _14__1_ d_lut_AOI21X1
ANOR2X1_19 [DC1.OUTPD_2_ _119__bF$buf4] _93_ d_lut_NOR2X1
AAOI21X1_9 [_107_ _119__bF$buf3 _93_] _14__2_ d_lut_AOI21X1
ANOR2X1_20 [DC1.OUTPD_3_ _119__bF$buf2] _94_ d_lut_NOR2X1
AAOI21X1_10 [_34_ _119__bF$buf1 _94_] _14__3_ d_lut_AOI21X1
ANOR2X1_21 [DC1.OUTPD_4_ _119__bF$buf0] _95_ d_lut_NOR2X1
AAOI21X1_11 [_40_ _119__bF$buf4 _95_] _14__4_ d_lut_AOI21X1
ANOR2X1_22 [DC1.OUTPD_5_ _119__bF$buf3] _96_ d_lut_NOR2X1
AAOI21X1_12 [_108_ _119__bF$buf2 _96_] _14__5_ d_lut_AOI21X1
ANOR2X1_23 [DC1.OUTPD_6_ _119__bF$buf1] _97_ d_lut_NOR2X1
AAOI21X1_13 [_112_ _119__bF$buf0 _97_] _14__6_ d_lut_AOI21X1
ANOR2X1_24 [DC1.OUTPD_7_ _119__bF$buf4] _98_ d_lut_NOR2X1
AAOI21X1_14 [_111_ _119__bF$buf3 _98_] _14__7_ d_lut_AOI21X1
AINVX1_13 [DC1.OUTPD_8_] _99_ d_lut_INVX1
ANOR2X1_25 [_99_ _119__bF$buf2] _14__8_ d_lut_NOR2X1
AINVX1_14 [DC1.OUTPD_9_] _100_ d_lut_INVX1
ANOR2X1_26 [_100_ _119__bF$buf1] _14__9_ d_lut_NOR2X1
AINVX1_15 [DC1.OUTPD_10_] _101_ d_lut_INVX1
ANOR2X1_27 [_101_ _119__bF$buf0] _14__10_ d_lut_NOR2X1
AINVX1_16 [DC1.OUTPD_11_] _102_ d_lut_INVX1
ANOR2X1_28 [_102_ _119__bF$buf4] _14__11_ d_lut_NOR2X1
AINVX1_17 [DC1.OUTPD_12_] _103_ d_lut_INVX1
ANOR2X1_29 [_103_ _119__bF$buf3] _14__12_ d_lut_NOR2X1
AINVX1_18 [DC1.OUTPD_13_] _104_ d_lut_INVX1
ANOR2X1_30 [_104_ _119__bF$buf2] _14__13_ d_lut_NOR2X1
AINVX1_19 [DC1.OUTPD_14_] _105_ d_lut_INVX1
ANOR2X1_31 [_105_ _119__bF$buf1] _14__14_ d_lut_NOR2X1
AINVX1_20 [DC1.OUTPD_15_] _106_ d_lut_INVX1
ANOR2X1_32 [_106_ _119__bF$buf0] _14__15_ d_lut_NOR2X1
ADFFPOSX1_2 _14__0_ clk_bF$buf4 NULL NULL DC1.OUTPD_0_ NULL ddflop
ADFFPOSX1_3 _14__1_ clk_bF$buf3 NULL NULL DC1.OUTPD_1_ NULL ddflop
ADFFPOSX1_4 _14__2_ clk_bF$buf2 NULL NULL DC1.OUTPD_2_ NULL ddflop
ADFFPOSX1_5 _14__3_ clk_bF$buf1 NULL NULL DC1.OUTPD_3_ NULL ddflop
ADFFPOSX1_6 _14__4_ clk_bF$buf0 NULL NULL DC1.OUTPD_4_ NULL ddflop
ADFFPOSX1_7 _14__5_ clk_bF$buf5 NULL NULL DC1.OUTPD_5_ NULL ddflop
ADFFPOSX1_8 _14__6_ clk_bF$buf4 NULL NULL DC1.OUTPD_6_ NULL ddflop
ADFFPOSX1_9 _14__7_ clk_bF$buf3 NULL NULL DC1.OUTPD_7_ NULL ddflop
ADFFPOSX1_10 _14__8_ clk_bF$buf2 NULL NULL DC1.OUTPD_8_ NULL ddflop
ADFFPOSX1_11 _14__9_ clk_bF$buf1 NULL NULL DC1.OUTPD_9_ NULL ddflop
ADFFPOSX1_12 _14__10_ clk_bF$buf0 NULL NULL DC1.OUTPD_10_ NULL ddflop
ADFFPOSX1_13 _14__11_ clk_bF$buf5 NULL NULL DC1.OUTPD_11_ NULL ddflop
ADFFPOSX1_14 _14__12_ clk_bF$buf4 NULL NULL DC1.OUTPD_12_ NULL ddflop
ADFFPOSX1_15 _14__13_ clk_bF$buf3 NULL NULL DC1.OUTPD_13_ NULL ddflop
ADFFPOSX1_16 _14__14_ clk_bF$buf2 NULL NULL DC1.OUTPD_14_ NULL ddflop
ADFFPOSX1_17 _14__15_ clk_bF$buf1 NULL NULL DC1.OUTPD_15_ NULL ddflop
ADFFPOSX1_18 _16__0_ clk_bF$buf0 NULL NULL DC1.WDATA_0_ NULL ddflop
ADFFPOSX1_19 _16__1_ clk_bF$buf5 NULL NULL DC1.WDATA_1_ NULL ddflop
ADFFPOSX1_20 _16__2_ clk_bF$buf4 NULL NULL DC1.WDATA_2_ NULL ddflop
ADFFPOSX1_21 _16__3_ clk_bF$buf3 NULL NULL DC1.WDATA_3_ NULL ddflop
ADFFPOSX1_22 _16__4_ clk_bF$buf2 NULL NULL DC1.WDATA_4_ NULL ddflop
ADFFPOSX1_23 _16__5_ clk_bF$buf1 NULL NULL DC1.WDATA_5_ NULL ddflop
ADFFPOSX1_24 _16__6_ clk_bF$buf0 NULL NULL DC1.WDATA_6_ NULL ddflop
ADFFPOSX1_25 _16__7_ clk_bF$buf5 NULL NULL DC1.WDATA_7_ NULL ddflop
ADFFPOSX1_26 _13_ clk_bF$buf4 NULL NULL DC1.IR NULL ddflop
ADFFPOSX1_27 _15_ clk_bF$buf3 NULL NULL DC1.OW NULL ddflop
AXOR2X1_3 [DPC1.DP_0_ DPC1.DPOP] _128__0_ d_lut_XOR2X1
AINVX1_21 [DPC1.DP_0_] _146_ d_lut_INVX1
ANOR2X1_33 [DC1.SGN_bF$buf3 _146_] _147_ d_lut_NOR2X1
AINVX8_1 [DC1.SGN_bF$buf2] _148_ d_lut_INVX8
ANOR2X1_34 [DPC1.DP_0_ _148_] _149_ d_lut_NOR2X1
AOAI21X1_31 [_147_ _149_ DPC1.DPOP] _150_ d_lut_OAI21X1
AXNOR2X1_2 [_150_ DPC1.DP_1_] _128__1_ d_lut_XNOR2X1
AAND2X2_11 [DPC1.DP_0_ DPC1.DP_1_] _151_ d_lut_AND2X2
AOR2X2_2 [_151_ DC1.SGN_bF$buf1] _152_ d_lut_OR2X2
AOAI21X1_32 [DPC1.DP_0_ DPC1.DP_1_ DC1.SGN_bF$buf0] _153_ d_lut_OAI21X1
ANAND3X1_9 [DPC1.DPOP _153_ _152_] _154_ d_lut_NAND3X1
AXNOR2X1_3 [_154_ DPC1.DP_2_] _128__2_ d_lut_XNOR2X1
AINVX2_7 [DPC1.DP_3_] _155_ d_lut_INVX2
ANAND2X1_20 [DPC1.DP_2_ _151_] _156_ d_lut_NAND2X1
ANOR3X1_4 [DPC1.DP_0_ DPC1.DP_1_ DPC1.DP_2_] _157_ d_lut_NOR3X1
AOAI21X1_33 [_157_ _148_ DPC1.DPOP] _158_ d_lut_OAI21X1
AAOI21X1_15 [_148_ _156_ _158_] _159_ d_lut_AOI21X1
AXNOR2X1_4 [_159_ _155_] _128__3_ d_lut_XNOR2X1
ANAND3X1_10 [DC1.SGN_bF$buf5 _155_ _157_] _160_ d_lut_NAND3X1
AAND2X2_12 [DPC1.DP_2_ DPC1.DP_3_] _161_ d_lut_AND2X2
ANAND2X1_21 [_161_ _151_] _162_ d_lut_NAND2X1
AOAI21X1_34 [_162_ DC1.SGN_bF$buf4 _160_] _163_ d_lut_OAI21X1
ANAND2X1_22 [DPC1.DPOP _163_] _164_ d_lut_NAND2X1
AXNOR2X1_5 [_164_ DPC1.DP_4_] _128__4_ d_lut_XNOR2X1
AINVX1_22 [DPC1.DP_4_] _165_ d_lut_INVX1
AOAI21X1_35 [_162_ _165_ _148_] _166_ d_lut_OAI21X1
AINVX2_8 [DPC1.DPOP] _167_ d_lut_INVX2
ANAND3X1_11 [_155_ _165_ _157_] _168_ d_lut_NAND3X1
AAOI21X1_16 [DC1.SGN_bF$buf3 _168_ _167_] _169_ d_lut_AOI21X1
ANAND2X1_23 [_166_ _169_] _170_ d_lut_NAND2X1
AXNOR2X1_6 [_170_ DPC1.DP_5_] _128__5_ d_lut_XNOR2X1
AOAI21X1_36 [_168_ DPC1.DP_5_ DC1.SGN_bF$buf2] _171_ d_lut_OAI21X1
ANAND2X1_24 [DPC1.DP_4_ DPC1.DP_5_] _172_ d_lut_NAND2X1
ANOR2X1_35 [_172_ _162_] _173_ d_lut_NOR2X1
AINVX1_23 [_173_] _174_ d_lut_INVX1
AAOI21X1_17 [_148_ _174_ _167_] _175_ d_lut_AOI21X1
ANAND2X1_25 [_171_ _175_] _176_ d_lut_NAND2X1
AXNOR2X1_7 [_176_ DPC1.DP_6_] _128__6_ d_lut_XNOR2X1
ANOR3X1_5 [DPC1.DP_5_ DPC1.DP_6_ _168_] _177_ d_lut_NOR3X1
ANAND2X1_26 [DPC1.DP_6_ _173_] _178_ d_lut_NAND2X1
AAOI21X1_18 [_148_ _178_ _167_] _179_ d_lut_AOI21X1
AOAI21X1_37 [_148_ _177_ _179_] _180_ d_lut_OAI21X1
AXNOR2X1_8 [_180_ DPC1.DP_7_] _128__7_ d_lut_XNOR2X1
AINVX1_24 [DPC1.DP_7_] _181_ d_lut_INVX1
AAND2X2_13 [_177_ _181_] _182_ d_lut_AND2X2
ANAND2X1_27 [DPC1.DP_6_ DPC1.DP_7_] _183_ d_lut_NAND2X1
AOR2X2_3 [_172_ _183_] _184_ d_lut_OR2X2
ANOR2X1_36 [_162_ _184_] _185_ d_lut_NOR2X1
ANOR2X1_37 [DC1.SGN_bF$buf1 _185_] _186_ d_lut_NOR2X1
ANOR2X1_38 [_167_ _186_] _187_ d_lut_NOR2X1
AOAI21X1_38 [_182_ _148_ _187_] _188_ d_lut_OAI21X1
AXNOR2X1_9 [_188_ DPC1.DP_8_] _128__8_ d_lut_XNOR2X1
AINVX1_25 [DPC1.DP_8_] _189_ d_lut_INVX1
ANAND3X1_12 [_181_ _189_ _177_] _190_ d_lut_NAND3X1
AOAI21X1_39 [DC1.SGN_bF$buf0 DPC1.DP_8_ _187_] _191_ d_lut_OAI21X1
AAOI21X1_19 [DC1.SGN_bF$buf5 _190_ _191_] _192_ d_lut_AOI21X1
AXOR2X1_4 [_192_ DPC1.DP_9_] _128__9_ d_lut_XOR2X1
ANOR2X1_39 [DPC1.DP_9_ _190_] _193_ d_lut_NOR2X1
ANAND3X1_13 [DPC1.DP_8_ DPC1.DP_9_ _185_] _194_ d_lut_NAND3X1
AAOI21X1_20 [_148_ _194_ _167_] _195_ d_lut_AOI21X1
AOAI21X1_40 [_193_ _148_ _195_] _196_ d_lut_OAI21X1
AXNOR2X1_10 [_196_ DPC1.DP_10_] _128__10_ d_lut_XNOR2X1
ANOR3X1_6 [DPC1.DP_9_ DPC1.DP_10_ _190_] _197_ d_lut_NOR3X1
AINVX1_26 [DPC1.DP_10_] _198_ d_lut_INVX1
AOAI21X1_41 [_194_ _198_ _148_] _199_ d_lut_OAI21X1
AAND2X2_14 [_199_ DPC1.DPOP] _200_ d_lut_AND2X2
AOAI21X1_42 [_148_ _197_ _200_] _201_ d_lut_OAI21X1
AXNOR2X1_11 [_201_ DPC1.DP_11_] _128__11_ d_lut_XNOR2X1
AINVX2_9 [DPC1.DP_12_] _129_ d_lut_INVX2
AINVX1_27 [DPC1.DP_11_] _130_ d_lut_INVX1
AAOI21X1_21 [_130_ _197_ _148_] _131_ d_lut_AOI21X1
ANOR3X1_7 [_198_ _130_ _194_] _132_ d_lut_NOR3X1
AOAI21X1_43 [_132_ DC1.SGN_bF$buf4 DPC1.DPOP] _133_ d_lut_OAI21X1
ANOR2X1_40 [_133_ _131_] _134_ d_lut_NOR2X1
AXNOR2X1_12 [_134_ _129_] _128__12_ d_lut_XNOR2X1
AINVX1_28 [DPC1.DP_13_] _135_ d_lut_INVX1
ANAND2X1_28 [_148_ _129_] _136_ d_lut_NAND2X1
ANAND2X1_29 [DC1.SGN_bF$buf3 DPC1.DP_12_] _137_ d_lut_NAND2X1
ANAND2X1_30 [_137_ _136_] _138_ d_lut_NAND2X1
ANOR3X1_8 [_133_ _138_ _131_] _139_ d_lut_NOR3X1
AXNOR2X1_13 [_139_ _135_] _128__13_ d_lut_XNOR2X1
AOAI21X1_44 [DC1.SGN_bF$buf2 DPC1.DP_13_ _137_] _140_ d_lut_OAI21X1
AAOI21X1_22 [DC1.SGN_bF$buf1 DPC1.DP_13_ _140_] _141_ d_lut_AOI21X1
ANAND3X1_14 [DPC1.DPOP _136_ _141_] _142_ d_lut_NAND3X1
AINVX1_29 [_142_] _143_ d_lut_INVX1
AOAI21X1_45 [_132_ DC1.SGN_bF$buf0 _143_] _144_ d_lut_OAI21X1
ANOR2X1_41 [_144_ _131_] _145_ d_lut_NOR2X1
AXOR2X1_5 [_145_ DPC1.DP_14_] _128__14_ d_lut_XOR2X1
ADFFPOSX1_28 _128__0_ clk_bF$buf2 NULL NULL DPC1.DP_0_ NULL ddflop
ADFFPOSX1_29 _128__1_ clk_bF$buf1 NULL NULL DPC1.DP_1_ NULL ddflop
ADFFPOSX1_30 _128__2_ clk_bF$buf0 NULL NULL DPC1.DP_2_ NULL ddflop
ADFFPOSX1_31 _128__3_ clk_bF$buf5 NULL NULL DPC1.DP_3_ NULL ddflop
ADFFPOSX1_32 _128__4_ clk_bF$buf4 NULL NULL DPC1.DP_4_ NULL ddflop
ADFFPOSX1_33 _128__5_ clk_bF$buf3 NULL NULL DPC1.DP_5_ NULL ddflop
ADFFPOSX1_34 _128__6_ clk_bF$buf2 NULL NULL DPC1.DP_6_ NULL ddflop
ADFFPOSX1_35 _128__7_ clk_bF$buf1 NULL NULL DPC1.DP_7_ NULL ddflop
ADFFPOSX1_36 _128__8_ clk_bF$buf0 NULL NULL DPC1.DP_8_ NULL ddflop
ADFFPOSX1_37 _128__9_ clk_bF$buf5 NULL NULL DPC1.DP_9_ NULL ddflop
ADFFPOSX1_38 _128__10_ clk_bF$buf4 NULL NULL DPC1.DP_10_ NULL ddflop
ADFFPOSX1_39 _128__11_ clk_bF$buf3 NULL NULL DPC1.DP_11_ NULL ddflop
ADFFPOSX1_40 _128__12_ clk_bF$buf2 NULL NULL DPC1.DP_12_ NULL ddflop
ADFFPOSX1_41 _128__13_ clk_bF$buf1 NULL NULL DPC1.DP_13_ NULL ddflop
ADFFPOSX1_42 _128__14_ clk_bF$buf0 NULL NULL DPC1.DP_14_ NULL ddflop
AAND2X2_15 [OPC1.INST_2_ OPC1.INST_1_] _212_ d_lut_AND2X2
AINVX2_10 [OPC1.INST_3_] _213_ d_lut_INVX2
AOAI21X1_46 [OPC1.INST_2_ OPC1.INST_1_ _213_] _214_ d_lut_OAI21X1
ANOR2X1_42 [_212_ _214_] _215_ d_lut_NOR2X1
ANAND2X1_31 [NEXTOP_2_ NEXTOP_1_] _216_ d_lut_NAND2X1
AINVX1_30 [_216_] _217_ d_lut_INVX1
ANOR2X1_43 [NEXTOP_2_ NEXTOP_1_] _218_ d_lut_NOR2X1
ANOR2X1_44 [_218_ _217_] _219_ d_lut_NOR2X1
AINVX1_31 [_219_] _220_ d_lut_INVX1
AOAI21X1_47 [_220_ NEXTOP_0_ _215_] _221_ d_lut_OAI21X1
AINVX1_32 [OPC1.INST_2_] _222_ d_lut_INVX1
ANAND2X1_32 [OPC1.INST_3_ _222_] _223_ d_lut_NAND2X1
ANOR2X1_45 [OPC1.INST_3_ DC1.SGN_bF$buf5] _224_ d_lut_NOR2X1
ANAND2X1_33 [_224_ _212_] _225_ d_lut_NAND2X1
AINVX2_11 [DC1.SGN_bF$buf4] _226_ d_lut_INVX2
AINVX4_3 [OPC1.INST_1_] _227_ d_lut_INVX4
ANAND3X1_15 [RF _226_ _227_] _228_ d_lut_NAND3X1
AINVX4_4 [DC1.IZ] _229_ d_lut_INVX4
ANAND2X1_34 [NEXTOP_0_ _229_] _230_ d_lut_NAND2X1
AOAI22X1_2 [_223_ _228_ _225_ _230_] _231_ d_lut_OAI22X1
ANAND2X1_35 [DC1.SGN_bF$buf3 _227_] _232_ d_lut_NAND2X1
AINVX2_12 [WF] _233_ d_lut_INVX2
ANOR2X1_46 [NEXTOP_0_ _233_] _234_ d_lut_NOR2X1
ANOR3X1_9 [_232_ _223_ _234_] _235_ d_lut_NOR3X1
AINVX1_33 [NEXTOP_2_] _236_ d_lut_INVX1
AINVX2_13 [NEXTOP_1_] _237_ d_lut_INVX2
AOAI21X1_48 [_236_ NEXTOP_0_ _237_] _238_ d_lut_OAI21X1
ANOR2X1_47 [OPC1.INST_3_ OPC1.INST_2_] _239_ d_lut_NOR2X1
ANAND3X1_16 [NEXTOP_0_ _227_ _239_] _240_ d_lut_NAND3X1
ANOR2X1_48 [_238_ _240_] _241_ d_lut_NOR2X1
ANOR3X1_10 [_241_ _235_ _231_] _242_ d_lut_NOR3X1
ANOR3X1_11 [NEXTOP_0_ OPC1.bracketcount_7_ _216_] _243_ d_lut_NOR3X1
ANAND2X1_36 [DC1.SGN_bF$buf2 OPC1.INST_1_] _244_ d_lut_NAND2X1
ANAND2X1_37 [OPC1.INST_3_ OPC1.INST_2_] _245_ d_lut_NAND2X1
AOR2X2_4 [_244_ _245_] _246_ d_lut_OR2X2
ANOR2X1_49 [_243_ _246_] _247_ d_lut_NOR2X1
AAND2X2_16 [OPC1.INST_3_ OPC1.INST_2_] _248_ d_lut_AND2X2
ANAND3X1_17 [DC1.SGN_bF$buf1 _227_ _248_] _249_ d_lut_NAND3X1
ANAND3X1_18 [_213_ DC1.SGN_bF$buf0 _212_] _250_ d_lut_NAND3X1
ANOR2X1_50 [NEXTOP_0_ _229_] _251_ d_lut_NOR2X1
AOAI21X1_49 [_250_ _251_ _249_] _252_ d_lut_OAI21X1
AINVX1_34 [NEXTOP_0_] _253_ d_lut_INVX1
ANAND3X1_19 [OPC1.INST_3_ OPC1.INST_1_ _222_] _254_ d_lut_NAND3X1
ANOR2X1_51 [_253_ _254_] _255_ d_lut_NOR2X1
ANOR3X1_12 [_247_ _255_ _252_] _256_ d_lut_NOR3X1
ANAND3X1_20 [_221_ _242_ _256_] OPC1.NEXTSTATE_0_ d_lut_NAND3X1
ANAND2X1_38 [OPC1.INST_2_ _213_] _257_ d_lut_NAND2X1
AOAI21X1_50 [_257_ _244_ _254_] _258_ d_lut_OAI21X1
ANOR3X1_13 [_232_ _233_ _223_] _259_ d_lut_NOR3X1
AOAI21X1_51 [_259_ _258_ NEXTOP_1_] _260_ d_lut_OAI21X1
ANAND2X1_39 [OPC1.INST_3_ _212_] _261_ d_lut_NAND2X1
AINVX1_35 [_261_] _262_ d_lut_INVX1
AAOI21X1_23 [_237_ _229_ _225_] _263_ d_lut_AOI21X1
ANOR2X1_52 [_262_ _263_] _264_ d_lut_NOR2X1
ANOR2X1_53 [_223_ _228_] _265_ d_lut_NOR2X1
ANOR3X1_14 [DC1.IZ _244_ _257_] _266_ d_lut_NOR3X1
ANAND2X1_40 [NEXTOP_1_ _236_] _267_ d_lut_NAND2X1
ANOR3X1_15 [_267_ _212_ _214_] _268_ d_lut_NOR3X1
ANOR3X1_16 [_266_ _265_ _268_] _269_ d_lut_NOR3X1
ANAND3X1_21 [_264_ _260_ _269_] OPC1.NEXTSTATE_1_ d_lut_NAND3X1
ANAND3X1_22 [NEXTOP_2_ NEXTOP_1_ NEXTOP_0_] _270_ d_lut_NAND3X1
AOAI21X1_52 [_270_ OPC1.bracketcount_7_ _226_] _271_ d_lut_OAI21X1
AOAI21X1_53 [_243_ _226_ _271_] _272_ d_lut_OAI21X1
ANAND2X1_41 [_262_ _272_] _273_ d_lut_NAND2X1
AOAI21X1_54 [_227_ _223_ _225_] _274_ d_lut_OAI21X1
AOAI21X1_55 [_259_ _274_ NEXTOP_2_] _275_ d_lut_OAI21X1
ANOR2X1_54 [NEXTOP_2_ _237_] _276_ d_lut_NOR2X1
ANOR3X1_17 [_214_ _212_ _276_] _277_ d_lut_NOR3X1
ANOR2X1_55 [NEXTOP_2_ _229_] _278_ d_lut_NOR2X1
ANOR3X1_18 [_244_ _257_ _278_] _279_ d_lut_NOR3X1
ANAND2X1_42 [_227_ _239_] _280_ d_lut_NAND2X1
AOAI22X1_3 [_280_ _218_ _225_ _229_] _281_ d_lut_OAI22X1
ANOR3X1_19 [_277_ _279_ _281_] _282_ d_lut_NOR3X1
ANAND3X1_23 [_273_ _275_ _282_] OPC1.NEXTSTATE_2_ d_lut_NAND3X1
AOAI21X1_56 [_217_ _218_ _215_] _283_ d_lut_OAI21X1
ANOR2X1_56 [_232_ _223_] _284_ d_lut_NOR2X1
ANAND2X1_43 [OPC1.INST_3_ _227_] _285_ d_lut_NAND2X1
AOAI21X1_57 [_285_ DC1.SGN_bF$buf5 _245_] _286_ d_lut_OAI21X1
AAOI21X1_24 [_233_ _284_ _286_] _287_ d_lut_AOI21X1
ANOR2X1_57 [_229_ _225_] _288_ d_lut_NOR2X1
AAOI21X1_25 [NEXTOP_2_ _253_ NEXTOP_1_] _289_ d_lut_AOI21X1
ANOR2X1_58 [_289_ _280_] _203_ d_lut_NOR2X1
ANOR3X1_20 [_203_ _266_ _288_] _204_ d_lut_NOR3X1
ANAND3X1_24 [_283_ _287_ _204_] OPC1.NEXTSTATE_3_ d_lut_NAND3X1
ANAND2X1_44 [_219_ _215_] _205_ d_lut_NAND2X1
ANOR2X1_59 [DC1.IZ _225_] _206_ d_lut_NOR2X1
AINVX1_36 [_250_] _207_ d_lut_INVX1
AAOI21X1_26 [DC1.IZ _207_ _206_] _208_ d_lut_AOI21X1
AOAI22X1_4 [_213_ _227_ _280_ _238_] _209_ d_lut_OAI22X1
ANOR2X1_60 [_259_ _209_] _210_ d_lut_NOR2X1
ANAND3X1_25 [_205_ _210_ _208_] OPC1.PCDELTA_0_ d_lut_NAND3X1
AINVX1_37 [_266_] _211_ d_lut_INVX1
AOAI21X1_58 [_243_ _246_ _211_] OPC1.PCDELTA_15_ d_lut_OAI21X1
AOAI21X1_59 [_229_ _225_ _211_] _202_ d_lut_OAI21X1
ADFFPOSX1_43 OPC1.NEXTSTATE_0_ clk_bF$buf5 NULL NULL DC1.SGN NULL ddflop
ADFFPOSX1_44 OPC1.NEXTSTATE_1_ clk_bF$buf4 NULL NULL OPC1.INST_1_ NULL ddflop
ADFFPOSX1_45 OPC1.NEXTSTATE_2_ clk_bF$buf3 NULL NULL OPC1.INST_2_ NULL ddflop
ADFFPOSX1_46 OPC1.NEXTSTATE_3_ clk_bF$buf2 NULL NULL OPC1.INST_3_ NULL ddflop
ABUFX2_61 [DC1.SGN_bF$buf4] OPC1.INST_0_ d_lut_BUFX2
ABUFX2_62 [OPC1.PCDELTA_15_bF$buf4] OPC1.PCDELTA_1_ d_lut_BUFX2
ABUFX2_63 [OPC1.PCDELTA_15_bF$buf3] OPC1.PCDELTA_2_ d_lut_BUFX2
ABUFX2_64 [OPC1.PCDELTA_15_bF$buf2] OPC1.PCDELTA_3_ d_lut_BUFX2
ABUFX2_65 [OPC1.PCDELTA_15_bF$buf1] OPC1.PCDELTA_4_ d_lut_BUFX2
ABUFX2_66 [OPC1.PCDELTA_15_bF$buf0] OPC1.PCDELTA_5_ d_lut_BUFX2
ABUFX2_67 [OPC1.PCDELTA_15_bF$buf4] OPC1.PCDELTA_6_ d_lut_BUFX2
ABUFX2_68 [OPC1.PCDELTA_15_bF$buf3] OPC1.PCDELTA_7_ d_lut_BUFX2
ABUFX2_69 [OPC1.PCDELTA_15_bF$buf2] OPC1.PCDELTA_8_ d_lut_BUFX2
ABUFX2_70 [OPC1.PCDELTA_15_bF$buf1] OPC1.PCDELTA_9_ d_lut_BUFX2
ABUFX2_71 [OPC1.PCDELTA_15_bF$buf0] OPC1.PCDELTA_10_ d_lut_BUFX2
ABUFX2_72 [OPC1.PCDELTA_15_bF$buf4] OPC1.PCDELTA_11_ d_lut_BUFX2
ABUFX2_73 [OPC1.PCDELTA_15_bF$buf3] OPC1.PCDELTA_12_ d_lut_BUFX2
ABUFX2_74 [OPC1.PCDELTA_15_bF$buf2] OPC1.PCDELTA_13_ d_lut_BUFX2
ABUFX2_75 [OPC1.PCDELTA_15_bF$buf1] OPC1.PCDELTA_14_ d_lut_BUFX2

.model todig_1v8 adc_bridge(in_high=1.2 in_low=0.6 rise_delay=10n fall_delay=10n)
.model toana_1v8 dac_bridge(out_high=1.8 out_low=0)

.model ddflop d_dff(ic=0 rise_delay=1n fall_delay=1n)
.model dzero d_pulldown(load=1p)
.model done d_pullup(load=1p)

AA2D1 [a_vdd] [vdd] todig_1v8
AA2D2 [a_clk] [clk] todig_1v8
AA2D3 [a_INPD_0_] [INPD_0_] todig_1v8
AA2D4 [a_INPD_1_] [INPD_1_] todig_1v8
AA2D5 [a_INPD_2_] [INPD_2_] todig_1v8
AA2D6 [a_INPD_3_] [INPD_3_] todig_1v8
AA2D7 [a_INPD_4_] [INPD_4_] todig_1v8
AA2D8 [a_INPD_5_] [INPD_5_] todig_1v8
AA2D9 [a_INPD_6_] [INPD_6_] todig_1v8
AA2D10 [a_INPD_7_] [INPD_7_] todig_1v8
AA2D11 [a_RDATA_0_] [RDATA_0_] todig_1v8
AA2D12 [a_RDATA_1_] [RDATA_1_] todig_1v8
AA2D13 [a_RDATA_2_] [RDATA_2_] todig_1v8
AA2D14 [a_RDATA_3_] [RDATA_3_] todig_1v8
AA2D15 [a_RDATA_4_] [RDATA_4_] todig_1v8
AA2D16 [a_RDATA_5_] [RDATA_5_] todig_1v8
AA2D17 [a_RDATA_6_] [RDATA_6_] todig_1v8
AA2D18 [a_RDATA_7_] [RDATA_7_] todig_1v8
AA2D19 [a_RF] [RF] todig_1v8
AA2D20 [a_WF] [WF] todig_1v8
AA2D21 [a_NEXTOP_0_] [NEXTOP_0_] todig_1v8
AA2D22 [a_NEXTOP_1_] [NEXTOP_1_] todig_1v8
AA2D23 [a_NEXTOP_2_] [NEXTOP_2_] todig_1v8
AD2A1 [IR] [a_IR] toana_1v8
AD2A2 [OW] [a_OW] toana_1v8
AD2A3 [OUTPD_0_] [a_OUTPD_0_] toana_1v8
AD2A4 [OUTPD_1_] [a_OUTPD_1_] toana_1v8
AD2A5 [OUTPD_2_] [a_OUTPD_2_] toana_1v8
AD2A6 [OUTPD_3_] [a_OUTPD_3_] toana_1v8
AD2A7 [OUTPD_4_] [a_OUTPD_4_] toana_1v8
AD2A8 [OUTPD_5_] [a_OUTPD_5_] toana_1v8
AD2A9 [OUTPD_6_] [a_OUTPD_6_] toana_1v8
AD2A10 [OUTPD_7_] [a_OUTPD_7_] toana_1v8
AD2A11 [OUTPD_8_] [a_OUTPD_8_] toana_1v8
AD2A12 [OUTPD_9_] [a_OUTPD_9_] toana_1v8
AD2A13 [OUTPD_10_] [a_OUTPD_10_] toana_1v8
AD2A14 [OUTPD_11_] [a_OUTPD_11_] toana_1v8
AD2A15 [OUTPD_12_] [a_OUTPD_12_] toana_1v8
AD2A16 [OUTPD_13_] [a_OUTPD_13_] toana_1v8
AD2A17 [OUTPD_14_] [a_OUTPD_14_] toana_1v8
AD2A18 [OUTPD_15_] [a_OUTPD_15_] toana_1v8
AD2A19 [reset] [a_reset] toana_1v8
AD2A20 [RD] [a_RD] toana_1v8
AD2A21 [WD] [a_WD] toana_1v8
AD2A22 [WDATA_0_] [a_WDATA_0_] toana_1v8
AD2A23 [WDATA_1_] [a_WDATA_1_] toana_1v8
AD2A24 [WDATA_2_] [a_WDATA_2_] toana_1v8
AD2A25 [WDATA_3_] [a_WDATA_3_] toana_1v8
AD2A26 [WDATA_4_] [a_WDATA_4_] toana_1v8
AD2A27 [WDATA_5_] [a_WDATA_5_] toana_1v8
AD2A28 [WDATA_6_] [a_WDATA_6_] toana_1v8
AD2A29 [WDATA_7_] [a_WDATA_7_] toana_1v8
AD2A30 [DP_0_] [a_DP_0_] toana_1v8
AD2A31 [DP_1_] [a_DP_1_] toana_1v8
AD2A32 [DP_2_] [a_DP_2_] toana_1v8
AD2A33 [DP_3_] [a_DP_3_] toana_1v8
AD2A34 [DP_4_] [a_DP_4_] toana_1v8
AD2A35 [DP_5_] [a_DP_5_] toana_1v8
AD2A36 [DP_6_] [a_DP_6_] toana_1v8
AD2A37 [DP_7_] [a_DP_7_] toana_1v8
AD2A38 [DP_8_] [a_DP_8_] toana_1v8
AD2A39 [DP_9_] [a_DP_9_] toana_1v8
AD2A40 [DP_10_] [a_DP_10_] toana_1v8
AD2A41 [DP_11_] [a_DP_11_] toana_1v8
AD2A42 [DP_12_] [a_DP_12_] toana_1v8
AD2A43 [DP_13_] [a_DP_13_] toana_1v8
AD2A44 [DP_14_] [a_DP_14_] toana_1v8
AD2A45 [PCDELTA_0_] [a_PCDELTA_0_] toana_1v8
AD2A46 [PCDELTA_1_] [a_PCDELTA_1_] toana_1v8
AD2A47 [PCDELTA_2_] [a_PCDELTA_2_] toana_1v8
AD2A48 [PCDELTA_3_] [a_PCDELTA_3_] toana_1v8
AD2A49 [PCDELTA_4_] [a_PCDELTA_4_] toana_1v8
AD2A50 [PCDELTA_5_] [a_PCDELTA_5_] toana_1v8
AD2A51 [PCDELTA_6_] [a_PCDELTA_6_] toana_1v8
AD2A52 [PCDELTA_7_] [a_PCDELTA_7_] toana_1v8
AD2A53 [PCDELTA_8_] [a_PCDELTA_8_] toana_1v8
AD2A54 [PCDELTA_9_] [a_PCDELTA_9_] toana_1v8
AD2A55 [PCDELTA_10_] [a_PCDELTA_10_] toana_1v8
AD2A56 [PCDELTA_11_] [a_PCDELTA_11_] toana_1v8
AD2A57 [PCDELTA_12_] [a_PCDELTA_12_] toana_1v8
AD2A58 [PCDELTA_13_] [a_PCDELTA_13_] toana_1v8
AD2A59 [PCDELTA_14_] [a_PCDELTA_14_] toana_1v8
AD2A60 [PCDELTA_15_] [a_PCDELTA_15_] toana_1v8

.ends BFCPU
 

* BUFX4 A
.model d_lut_BUFX4 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "01")
* INVX1 (!A)
.model d_lut_INVX1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "10")
* NAND2X1 (!(A B))
.model d_lut_NAND2X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "1110")
* OR2X2 (A+B)
.model d_lut_OR2X2 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "0111")
* NOR2X1 (!(A+B))
.model d_lut_NOR2X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "1000")
* AND2X2 (A B)
.model d_lut_AND2X2 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "0001")
* BUFX2 A
.model d_lut_BUFX2 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "01")
* DFFPOSX1 DS0000
* INVX4 (!A)
.model d_lut_INVX4 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "10")
* INVX2 (!A)
.model d_lut_INVX2 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "10")
* NAND3X1 (!((A B) C))
.model d_lut_NAND3X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "11111110")
* XOR2X1 (A^B)
.model d_lut_XOR2X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "0110")
* OAI21X1 (!((A+B) C))
.model d_lut_OAI21X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "11111000")
* AOI22X1 (!((A B)+(C D)))
.model d_lut_AOI22X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "1110111011100000")
* XNOR2X1 (!(A^B))
.model d_lut_XNOR2X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "1001")
* MUX2X1 (!((S A) + (!S B)))
.model d_lut_MUX2X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "11001010")
* OAI22X1 (!((A+B) (C+D)))
.model d_lut_OAI22X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "1111100010001000")
* NOR3X1 (!((A+B)+C))
.model d_lut_NOR3X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "10000000")
* AOI21X1 (!((A B)+C))
.model d_lut_AOI21X1 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "11100000")
* INVX8 (!A)
.model d_lut_INVX8 d_lut (rise_delay=1n fall_delay=1n input_load=10f
+ table_values "10")
.end
