magic
tech scmos
timestamp 1537539148
<< metal1 >>
rect 476 1203 477 1207
rect 481 1203 482 1207
rect 486 1203 488 1207
rect 462 1188 478 1191
rect 94 1168 102 1171
rect 733 1168 734 1172
rect 1078 1166 1082 1168
rect 1102 1168 1110 1171
rect 1102 1166 1106 1168
rect 1150 1166 1154 1168
rect 1206 1166 1210 1168
rect 1222 1168 1234 1171
rect 1222 1162 1225 1168
rect 1230 1166 1234 1168
rect 1270 1166 1274 1168
rect 502 1158 510 1161
rect 118 1148 129 1151
rect 286 1148 297 1151
rect 118 1142 121 1148
rect 286 1142 289 1148
rect 578 1148 585 1151
rect 734 1148 750 1151
rect 814 1148 825 1151
rect 242 1138 249 1141
rect 638 1141 641 1148
rect 814 1142 817 1148
rect 934 1148 942 1151
rect 1298 1148 1305 1151
rect 630 1138 641 1141
rect 958 1138 977 1141
rect 1010 1138 1025 1141
rect 1030 1138 1049 1141
rect 1082 1138 1089 1141
rect 1166 1138 1185 1141
rect 1250 1138 1254 1141
rect 110 1128 121 1131
rect 262 1128 281 1131
rect 598 1131 602 1136
rect 586 1128 602 1131
rect 942 1128 945 1138
rect 990 1128 1014 1131
rect 1074 1118 1075 1122
rect 1098 1118 1099 1122
rect 1122 1118 1123 1122
rect 1146 1118 1147 1122
rect 1213 1118 1214 1122
rect 1237 1118 1238 1122
rect 1462 1118 1486 1121
rect 988 1103 989 1107
rect 993 1103 994 1107
rect 998 1103 1000 1107
rect 1058 1088 1059 1092
rect 110 1078 121 1081
rect 190 1078 201 1081
rect 138 1068 153 1071
rect 430 1071 433 1081
rect 558 1078 577 1081
rect 414 1068 433 1071
rect 446 1068 486 1071
rect 614 1071 617 1081
rect 654 1078 673 1081
rect 678 1078 690 1081
rect 686 1077 690 1078
rect 1118 1072 1121 1081
rect 598 1068 617 1071
rect 634 1068 641 1071
rect 942 1068 950 1071
rect 990 1068 1001 1071
rect 38 1058 46 1061
rect 118 1061 121 1068
rect 118 1058 129 1061
rect 134 1058 137 1068
rect 246 1058 254 1061
rect 342 1058 358 1061
rect 426 1058 433 1061
rect 502 1058 521 1061
rect 934 1058 942 1061
rect 990 1061 993 1068
rect 974 1058 993 1061
rect 1082 1058 1097 1061
rect 1210 1058 1222 1061
rect 1458 1058 1465 1061
rect 614 1051 617 1058
rect 614 1048 625 1051
rect 1098 1048 1102 1052
rect 933 1038 934 1042
rect 181 1018 182 1022
rect 794 1018 795 1022
rect 1197 1018 1198 1022
rect 476 1003 477 1007
rect 481 1003 482 1007
rect 486 1003 488 1007
rect 1140 968 1142 972
rect 990 958 998 961
rect 118 941 121 948
rect 134 942 137 951
rect 226 948 233 951
rect 446 948 454 951
rect 118 938 129 941
rect 446 941 449 948
rect 738 948 745 951
rect 822 948 830 951
rect 970 948 977 951
rect 1070 948 1086 951
rect 138 938 153 941
rect 446 938 465 941
rect 550 938 558 941
rect 766 938 777 941
rect 958 938 969 941
rect 1078 938 1097 941
rect 94 931 98 933
rect 382 931 386 933
rect 1078 932 1081 938
rect 94 928 105 931
rect 110 928 121 931
rect 382 928 390 931
rect 406 928 417 931
rect 438 928 446 931
rect 694 928 713 931
rect 990 918 998 921
rect 988 903 989 907
rect 993 903 994 907
rect 998 903 1000 907
rect 94 878 105 881
rect 110 878 121 881
rect 246 878 257 881
rect 294 878 305 881
rect 646 878 657 881
rect 662 878 681 881
rect 94 877 98 878
rect 646 877 650 878
rect 310 868 322 871
rect 502 868 534 871
rect 694 868 702 871
rect 118 861 121 868
rect 118 858 129 861
rect 254 861 257 868
rect 254 858 265 861
rect 270 858 278 861
rect 294 861 297 868
rect 286 858 297 861
rect 310 862 313 868
rect 702 858 721 861
rect 758 861 761 871
rect 854 868 873 871
rect 898 868 905 871
rect 1086 862 1089 871
rect 750 858 761 861
rect 790 858 810 861
rect 986 858 1009 861
rect 1126 861 1129 871
rect 1118 858 1129 861
rect 1150 858 1169 861
rect 1434 858 1441 861
rect 806 856 810 858
rect 806 848 817 851
rect 1150 848 1153 858
rect 814 842 817 848
rect 942 838 950 841
rect 476 803 477 807
rect 481 803 482 807
rect 486 803 488 807
rect 546 768 547 772
rect 454 758 462 761
rect 154 748 161 751
rect 254 748 262 751
rect 494 748 510 751
rect 694 748 726 751
rect 842 748 846 751
rect 1030 748 1041 751
rect 166 738 185 741
rect 514 738 521 741
rect 670 741 673 748
rect 670 738 684 741
rect 814 738 825 741
rect 1038 738 1041 748
rect 1062 738 1065 748
rect 1178 748 1185 751
rect 1250 748 1257 751
rect 1450 748 1457 751
rect 182 728 185 738
rect 422 731 425 738
rect 822 732 825 738
rect 422 728 436 731
rect 122 718 124 722
rect 982 718 990 721
rect 988 703 989 707
rect 993 703 994 707
rect 998 703 1000 707
rect 897 688 902 692
rect 70 678 86 681
rect 754 678 761 681
rect 802 678 817 681
rect 910 681 913 688
rect 910 678 934 681
rect 1126 678 1134 681
rect 1306 678 1322 681
rect 70 674 74 678
rect 142 668 154 671
rect 378 668 385 671
rect 434 668 441 671
rect 494 668 505 671
rect 622 668 649 671
rect 666 668 681 671
rect 690 668 697 671
rect 846 668 881 671
rect 1110 671 1113 678
rect 1318 674 1322 678
rect 1102 668 1113 671
rect 1182 668 1193 671
rect 1298 668 1299 672
rect 46 658 58 661
rect 250 658 273 661
rect 342 658 350 661
rect 502 661 505 668
rect 466 658 481 661
rect 502 658 513 661
rect 586 658 601 661
rect 702 658 721 661
rect 830 658 849 661
rect 1110 658 1121 661
rect 1162 658 1169 661
rect 1222 658 1238 661
rect 1334 658 1345 661
rect 1398 658 1414 661
rect 54 657 58 658
rect 718 648 721 658
rect 1334 657 1338 658
rect 922 648 929 651
rect 826 638 827 642
rect 1454 618 1462 621
rect 476 603 477 607
rect 481 603 482 607
rect 486 603 488 607
rect 341 588 342 592
rect 470 588 478 591
rect 501 588 502 592
rect 538 568 541 572
rect 875 568 878 572
rect 118 558 129 561
rect 302 558 313 561
rect 318 558 326 561
rect 398 558 409 561
rect 626 558 630 562
rect 690 558 694 562
rect 990 558 1006 561
rect 1236 558 1238 562
rect 118 552 121 558
rect 54 548 65 551
rect 318 548 337 551
rect 374 548 393 551
rect 446 548 454 551
rect 474 548 497 551
rect 54 542 57 548
rect 82 538 89 541
rect 198 538 217 541
rect 422 541 425 548
rect 630 548 638 551
rect 670 548 681 551
rect 1102 548 1113 551
rect 1350 551 1354 553
rect 422 538 433 541
rect 638 538 646 541
rect 678 538 681 548
rect 858 538 859 542
rect 950 538 966 541
rect 1102 538 1105 548
rect 1174 538 1177 548
rect 1350 548 1361 551
rect 94 531 97 538
rect 94 528 110 531
rect 230 528 249 531
rect 414 528 417 538
rect 950 528 953 538
rect 1150 528 1161 531
rect 1334 531 1338 536
rect 1322 528 1338 531
rect 1158 522 1161 528
rect 394 518 395 522
rect 1093 518 1094 522
rect 988 503 989 507
rect 993 503 994 507
rect 998 503 1000 507
rect 182 488 190 491
rect 474 488 475 492
rect 1018 488 1020 492
rect 134 468 153 471
rect 398 471 401 481
rect 442 478 446 482
rect 498 478 505 481
rect 398 468 406 471
rect 550 468 569 471
rect 614 468 634 471
rect 742 468 750 471
rect 918 471 922 474
rect 918 468 929 471
rect 994 468 1001 471
rect 1082 468 1097 471
rect 1278 468 1286 471
rect 38 458 46 461
rect 254 458 262 461
rect 374 458 382 461
rect 814 458 822 461
rect 1130 458 1145 461
rect 1290 458 1297 461
rect 94 451 98 454
rect 94 448 105 451
rect 250 448 254 452
rect 478 448 505 451
rect 946 448 948 452
rect 1142 448 1145 458
rect 1250 448 1254 452
rect 182 438 198 441
rect 222 438 242 441
rect 1222 438 1242 441
rect 222 428 225 438
rect 1222 428 1225 438
rect 476 403 477 407
rect 481 403 482 407
rect 486 403 488 407
rect 229 388 230 392
rect 818 388 820 392
rect 874 388 876 392
rect 98 368 105 371
rect 1018 368 1019 372
rect 130 358 137 361
rect 422 358 433 361
rect 1150 358 1161 361
rect 1202 358 1206 361
rect 38 348 81 351
rect 194 348 201 351
rect 218 348 225 351
rect 254 348 262 351
rect 446 348 454 351
rect 458 348 462 351
rect 46 338 70 341
rect 174 338 193 341
rect 374 341 377 348
rect 698 348 702 351
rect 730 348 737 351
rect 762 348 769 351
rect 990 348 1014 351
rect 1226 348 1233 351
rect 366 338 377 341
rect 630 338 642 341
rect 702 338 721 341
rect 990 341 993 348
rect 982 338 993 341
rect 1002 338 1009 341
rect 1126 338 1137 341
rect 1174 338 1193 341
rect 1302 338 1310 341
rect 630 332 633 338
rect 1206 332 1209 338
rect 66 328 73 331
rect 1206 328 1214 332
rect 149 318 150 322
rect 178 318 179 322
rect 329 318 342 321
rect 586 318 587 322
rect 1284 318 1286 322
rect 988 303 989 307
rect 993 303 994 307
rect 998 303 1000 307
rect 398 288 406 291
rect 982 288 990 291
rect 166 278 182 281
rect 578 278 588 281
rect 814 278 822 281
rect 918 278 929 281
rect 1154 278 1161 281
rect 1230 278 1238 281
rect 814 277 818 278
rect 94 271 98 274
rect 94 268 105 271
rect 150 268 161 271
rect 350 268 358 271
rect 366 268 377 271
rect 446 268 481 271
rect 830 268 841 271
rect 1226 268 1233 271
rect 214 258 233 261
rect 250 258 262 261
rect 310 261 313 268
rect 310 258 321 261
rect 378 258 385 261
rect 478 261 481 268
rect 478 258 497 261
rect 502 258 521 261
rect 534 258 566 261
rect 842 258 857 261
rect 994 258 1009 261
rect 1098 258 1110 261
rect 1126 258 1145 261
rect 1150 258 1169 261
rect 1234 258 1241 261
rect 1294 258 1305 261
rect 1470 258 1478 261
rect 518 248 521 258
rect 1126 248 1129 258
rect 1182 256 1186 258
rect 795 238 798 242
rect 1290 238 1291 242
rect 237 218 238 222
rect 1114 218 1115 222
rect 476 203 477 207
rect 481 203 482 207
rect 486 203 488 207
rect 362 188 363 192
rect 470 188 486 191
rect 541 188 542 192
rect 210 178 211 182
rect 450 168 465 171
rect 682 158 689 161
rect 982 158 1006 161
rect 1046 158 1057 161
rect 1066 158 1070 162
rect 558 152 562 154
rect 86 148 113 151
rect 118 148 145 151
rect 254 148 262 151
rect 290 148 294 151
rect 342 148 350 151
rect 366 148 374 151
rect 402 148 409 151
rect 418 148 433 151
rect 498 148 505 151
rect 634 148 649 151
rect 722 148 737 151
rect 1002 148 1017 151
rect 1070 148 1078 151
rect 1094 148 1126 151
rect 1162 148 1166 151
rect 1170 148 1177 151
rect 1334 148 1342 151
rect 86 142 89 148
rect 42 138 57 141
rect 310 138 329 141
rect 326 128 329 138
rect 1438 133 1442 138
rect 346 128 353 131
rect 738 128 745 131
rect 1114 128 1121 131
rect 882 118 883 122
rect 1284 118 1286 122
rect 1454 118 1470 121
rect 988 103 989 107
rect 993 103 994 107
rect 998 103 1000 107
rect 716 88 718 92
rect 869 88 870 92
rect 1074 88 1081 91
rect 54 78 62 81
rect 318 78 326 81
rect 490 78 497 81
rect 846 78 854 81
rect 98 68 105 71
rect 226 68 230 71
rect 278 68 289 71
rect 362 68 377 71
rect 394 68 409 71
rect 514 68 521 71
rect 542 68 569 71
rect 750 68 761 71
rect 818 68 825 71
rect 926 71 929 81
rect 998 78 1006 81
rect 926 68 934 71
rect 998 71 1001 78
rect 990 68 1001 71
rect 1018 68 1036 71
rect 1054 68 1062 71
rect 1134 68 1153 71
rect 1174 68 1185 71
rect 38 58 81 61
rect 86 58 94 61
rect 118 58 129 61
rect 182 58 198 61
rect 274 58 278 61
rect 314 58 329 61
rect 462 58 470 61
rect 510 58 526 61
rect 894 58 905 61
rect 1046 58 1054 61
rect 1094 58 1113 61
rect 1214 58 1230 61
rect 446 51 449 58
rect 438 48 449 51
rect 958 48 969 51
rect 286 38 294 41
rect 778 38 780 42
rect 946 38 947 42
rect 476 3 477 7
rect 481 3 482 7
rect 486 3 488 7
<< m2contact >>
rect 472 1203 476 1207
rect 477 1203 481 1207
rect 482 1203 486 1207
rect 158 1188 162 1192
rect 182 1188 186 1192
rect 230 1188 234 1192
rect 310 1188 314 1192
rect 334 1188 338 1192
rect 390 1188 394 1192
rect 414 1188 418 1192
rect 438 1188 442 1192
rect 478 1188 482 1192
rect 694 1188 698 1192
rect 1318 1188 1322 1192
rect 1342 1188 1346 1192
rect 1366 1188 1370 1192
rect 1390 1188 1394 1192
rect 1414 1188 1418 1192
rect 1438 1188 1442 1192
rect 206 1178 210 1182
rect 686 1178 690 1182
rect 102 1168 106 1172
rect 662 1168 666 1172
rect 734 1168 738 1172
rect 790 1168 794 1172
rect 1078 1168 1082 1172
rect 1110 1168 1114 1172
rect 1150 1168 1154 1172
rect 1206 1168 1210 1172
rect 1270 1168 1274 1172
rect 510 1158 514 1162
rect 638 1158 642 1162
rect 718 1158 722 1162
rect 774 1158 778 1162
rect 1126 1158 1130 1162
rect 1222 1158 1226 1162
rect 38 1148 42 1152
rect 134 1148 138 1152
rect 142 1148 146 1152
rect 166 1148 170 1152
rect 190 1148 194 1152
rect 214 1148 218 1152
rect 238 1148 242 1152
rect 270 1148 274 1152
rect 318 1148 322 1152
rect 366 1148 370 1152
rect 374 1148 378 1152
rect 398 1148 402 1152
rect 422 1148 426 1152
rect 446 1148 450 1152
rect 550 1147 554 1151
rect 574 1148 578 1152
rect 638 1148 642 1152
rect 646 1148 650 1152
rect 670 1148 674 1152
rect 710 1148 714 1152
rect 750 1148 754 1152
rect 758 1148 762 1152
rect 766 1148 770 1152
rect 782 1148 786 1152
rect 118 1138 122 1142
rect 238 1138 242 1142
rect 286 1138 290 1142
rect 486 1138 490 1142
rect 518 1138 522 1142
rect 622 1138 626 1142
rect 862 1147 866 1151
rect 942 1148 946 1152
rect 966 1148 970 1152
rect 982 1148 986 1152
rect 1038 1148 1042 1152
rect 1174 1148 1178 1152
rect 1294 1148 1298 1152
rect 1326 1148 1330 1152
rect 1350 1148 1354 1152
rect 1374 1148 1378 1152
rect 1398 1148 1402 1152
rect 1422 1148 1426 1152
rect 1446 1148 1450 1152
rect 742 1138 746 1142
rect 750 1138 754 1142
rect 790 1138 794 1142
rect 806 1138 810 1142
rect 814 1138 818 1142
rect 830 1138 834 1142
rect 846 1138 850 1142
rect 942 1138 946 1142
rect 1006 1138 1010 1142
rect 1062 1138 1066 1142
rect 1078 1138 1082 1142
rect 1110 1138 1114 1142
rect 1134 1138 1138 1142
rect 1222 1138 1226 1142
rect 1246 1138 1250 1142
rect 1254 1138 1258 1142
rect 30 1128 34 1132
rect 102 1128 106 1132
rect 286 1128 290 1132
rect 582 1128 586 1132
rect 950 1128 954 1132
rect 1014 1128 1018 1132
rect 1054 1128 1058 1132
rect 1158 1128 1162 1132
rect 1198 1128 1202 1132
rect 254 1118 258 1122
rect 350 1118 354 1122
rect 502 1118 506 1122
rect 614 1118 618 1122
rect 926 1118 930 1122
rect 1070 1118 1074 1122
rect 1094 1118 1098 1122
rect 1118 1118 1122 1122
rect 1142 1118 1146 1122
rect 1190 1118 1194 1122
rect 1214 1118 1218 1122
rect 1238 1118 1242 1122
rect 1270 1118 1274 1122
rect 1486 1118 1490 1122
rect 984 1103 988 1107
rect 989 1103 993 1107
rect 994 1103 998 1107
rect 94 1088 98 1092
rect 302 1088 306 1092
rect 398 1088 402 1092
rect 550 1088 554 1092
rect 686 1088 690 1092
rect 790 1088 794 1092
rect 894 1088 898 1092
rect 910 1088 914 1092
rect 1054 1088 1058 1092
rect 1294 1088 1298 1092
rect 1310 1088 1314 1092
rect 1374 1088 1378 1092
rect 1398 1088 1402 1092
rect 1414 1088 1418 1092
rect 1438 1088 1442 1092
rect 1478 1088 1482 1092
rect 30 1078 34 1082
rect 102 1078 106 1082
rect 206 1078 210 1082
rect 422 1078 426 1082
rect 118 1068 122 1072
rect 134 1068 138 1072
rect 222 1068 226 1072
rect 350 1068 354 1072
rect 510 1078 514 1082
rect 582 1078 586 1082
rect 606 1078 610 1082
rect 486 1068 490 1072
rect 542 1068 546 1072
rect 782 1078 786 1082
rect 806 1078 810 1082
rect 630 1068 634 1072
rect 766 1068 770 1072
rect 822 1068 826 1072
rect 862 1068 866 1072
rect 870 1068 874 1072
rect 902 1068 906 1072
rect 950 1068 954 1072
rect 1030 1068 1034 1072
rect 1086 1068 1090 1072
rect 1118 1068 1122 1072
rect 1206 1068 1210 1072
rect 1214 1068 1218 1072
rect 1230 1068 1234 1072
rect 1246 1068 1250 1072
rect 1262 1068 1266 1072
rect 46 1058 50 1062
rect 62 1058 66 1062
rect 166 1058 170 1062
rect 174 1058 178 1062
rect 254 1058 258 1062
rect 270 1058 274 1062
rect 358 1058 362 1062
rect 406 1058 410 1062
rect 422 1058 426 1062
rect 454 1058 458 1062
rect 526 1058 530 1062
rect 534 1058 538 1062
rect 566 1058 570 1062
rect 590 1058 594 1062
rect 614 1058 618 1062
rect 630 1058 634 1062
rect 662 1058 666 1062
rect 718 1058 722 1062
rect 742 1058 746 1062
rect 798 1058 802 1062
rect 830 1058 834 1062
rect 854 1058 858 1062
rect 878 1058 882 1062
rect 942 1058 946 1062
rect 958 1058 962 1062
rect 1006 1058 1010 1062
rect 1022 1058 1026 1062
rect 1038 1058 1042 1062
rect 1046 1058 1050 1062
rect 1070 1058 1074 1062
rect 1078 1058 1082 1062
rect 1134 1058 1138 1062
rect 1142 1058 1146 1062
rect 1166 1058 1170 1062
rect 1198 1058 1202 1062
rect 1206 1058 1210 1062
rect 1222 1058 1226 1062
rect 1254 1058 1258 1062
rect 1278 1058 1282 1062
rect 1326 1058 1330 1062
rect 1350 1058 1354 1062
rect 1358 1058 1362 1062
rect 1382 1058 1386 1062
rect 1430 1058 1434 1062
rect 1454 1058 1458 1062
rect 654 1048 658 1052
rect 838 1048 842 1052
rect 848 1048 852 1052
rect 894 1048 898 1052
rect 918 1048 922 1052
rect 1094 1048 1098 1052
rect 1110 1048 1114 1052
rect 1182 1048 1186 1052
rect 1238 1048 1242 1052
rect 1270 1048 1274 1052
rect 934 1038 938 1042
rect 182 1018 186 1022
rect 526 1018 530 1022
rect 790 1018 794 1022
rect 806 1018 810 1022
rect 1014 1018 1018 1022
rect 1126 1018 1130 1022
rect 1158 1018 1162 1022
rect 1198 1018 1202 1022
rect 472 1003 476 1007
rect 477 1003 481 1007
rect 482 1003 486 1007
rect 94 988 98 992
rect 262 988 266 992
rect 286 988 290 992
rect 382 988 386 992
rect 582 988 586 992
rect 926 988 930 992
rect 1030 988 1034 992
rect 1230 988 1234 992
rect 1294 988 1298 992
rect 1318 988 1322 992
rect 1358 988 1362 992
rect 1374 988 1378 992
rect 1398 988 1402 992
rect 390 968 394 972
rect 590 968 594 972
rect 1142 968 1146 972
rect 766 958 770 962
rect 798 958 802 962
rect 830 958 834 962
rect 958 958 962 962
rect 998 958 1002 962
rect 1222 958 1226 962
rect 38 948 42 952
rect 62 948 66 952
rect 118 948 122 952
rect 166 948 170 952
rect 198 947 202 951
rect 222 948 226 952
rect 270 948 274 952
rect 326 948 330 952
rect 350 948 354 952
rect 390 948 394 952
rect 454 948 458 952
rect 478 948 482 952
rect 526 948 530 952
rect 534 948 538 952
rect 566 948 570 952
rect 134 938 138 942
rect 654 947 658 951
rect 702 948 706 952
rect 734 948 738 952
rect 750 948 754 952
rect 782 948 786 952
rect 814 948 818 952
rect 830 948 834 952
rect 862 947 866 951
rect 942 948 946 952
rect 966 948 970 952
rect 1022 948 1026 952
rect 1046 948 1050 952
rect 1054 948 1058 952
rect 1062 948 1066 952
rect 1086 948 1090 952
rect 1102 948 1106 952
rect 1190 948 1194 952
rect 1206 948 1210 952
rect 1246 948 1250 952
rect 1254 948 1258 952
rect 1278 948 1282 952
rect 1310 948 1314 952
rect 1334 948 1338 952
rect 1342 948 1346 952
rect 1390 948 1394 952
rect 1414 948 1418 952
rect 1438 948 1442 952
rect 1462 948 1466 952
rect 518 938 522 942
rect 558 938 562 942
rect 638 938 642 942
rect 726 938 730 942
rect 742 938 746 942
rect 806 938 810 942
rect 846 938 850 942
rect 934 938 938 942
rect 1110 938 1114 942
rect 1158 938 1162 942
rect 1182 938 1186 942
rect 1198 938 1202 942
rect 30 928 34 932
rect 390 928 394 932
rect 422 928 426 932
rect 430 928 434 932
rect 446 928 450 932
rect 502 928 506 932
rect 686 928 690 932
rect 718 928 722 932
rect 1078 928 1082 932
rect 1086 928 1090 932
rect 1166 928 1170 932
rect 1238 928 1242 932
rect 150 918 154 922
rect 510 918 514 922
rect 798 918 802 922
rect 926 918 930 922
rect 998 918 1002 922
rect 1174 918 1178 922
rect 1222 918 1226 922
rect 1270 918 1274 922
rect 984 903 988 907
rect 989 903 993 907
rect 994 903 998 907
rect 94 888 98 892
rect 230 888 234 892
rect 406 888 410 892
rect 414 888 418 892
rect 646 888 650 892
rect 718 888 722 892
rect 782 888 786 892
rect 790 888 794 892
rect 846 888 850 892
rect 974 888 978 892
rect 1030 888 1034 892
rect 1390 888 1394 892
rect 1462 888 1466 892
rect 30 878 34 882
rect 238 878 242 882
rect 310 878 314 882
rect 686 878 690 882
rect 710 878 714 882
rect 838 878 842 882
rect 926 878 930 882
rect 118 868 122 872
rect 254 868 258 872
rect 294 868 298 872
rect 534 868 538 872
rect 566 868 570 872
rect 702 868 706 872
rect 726 868 730 872
rect 38 858 42 862
rect 134 858 138 862
rect 174 858 178 862
rect 198 858 202 862
rect 278 858 282 862
rect 310 858 314 862
rect 342 859 346 863
rect 374 858 378 862
rect 478 859 482 863
rect 550 858 554 862
rect 590 858 594 862
rect 670 858 674 862
rect 734 858 738 862
rect 798 868 802 872
rect 894 868 898 872
rect 966 868 970 872
rect 1022 868 1026 872
rect 1054 868 1058 872
rect 1062 868 1066 872
rect 1094 868 1098 872
rect 766 858 770 862
rect 814 858 818 862
rect 862 858 866 862
rect 886 858 890 862
rect 910 858 914 862
rect 950 858 954 862
rect 982 858 986 862
rect 1046 858 1050 862
rect 1070 858 1074 862
rect 1086 858 1090 862
rect 1102 858 1106 862
rect 1150 868 1154 872
rect 1182 868 1186 872
rect 1294 868 1298 872
rect 1134 858 1138 862
rect 1174 858 1178 862
rect 1214 859 1218 863
rect 1246 858 1250 862
rect 1310 859 1314 863
rect 1406 858 1410 862
rect 1430 858 1434 862
rect 1478 858 1482 862
rect 782 848 786 852
rect 870 848 874 852
rect 926 848 930 852
rect 958 848 962 852
rect 1086 848 1090 852
rect 1158 848 1162 852
rect 814 838 818 842
rect 822 838 826 842
rect 950 838 954 842
rect 1278 838 1282 842
rect 934 828 938 832
rect 814 818 818 822
rect 1030 818 1034 822
rect 1374 818 1378 822
rect 472 803 476 807
rect 477 803 481 807
rect 482 803 486 807
rect 230 788 234 792
rect 614 788 618 792
rect 646 788 650 792
rect 894 788 898 792
rect 942 788 946 792
rect 1166 788 1170 792
rect 1198 788 1202 792
rect 1398 788 1402 792
rect 1422 778 1426 782
rect 94 768 98 772
rect 438 768 442 772
rect 542 768 546 772
rect 582 768 586 772
rect 606 768 610 772
rect 638 768 642 772
rect 774 768 778 772
rect 814 768 818 772
rect 886 768 890 772
rect 902 768 906 772
rect 1222 768 1226 772
rect 462 758 466 762
rect 502 758 506 762
rect 558 758 562 762
rect 566 758 570 762
rect 622 758 626 762
rect 654 758 658 762
rect 742 758 746 762
rect 798 758 802 762
rect 830 758 834 762
rect 862 758 866 762
rect 870 758 874 762
rect 982 758 986 762
rect 1062 758 1066 762
rect 38 748 42 752
rect 62 748 66 752
rect 150 748 154 752
rect 206 748 210 752
rect 214 748 218 752
rect 262 748 266 752
rect 286 748 290 752
rect 374 747 378 751
rect 422 748 426 752
rect 446 748 450 752
rect 486 748 490 752
rect 510 748 514 752
rect 526 748 530 752
rect 542 748 546 752
rect 574 748 578 752
rect 590 748 594 752
rect 614 748 618 752
rect 646 748 650 752
rect 670 748 674 752
rect 726 748 730 752
rect 758 748 762 752
rect 822 748 826 752
rect 838 748 842 752
rect 846 748 850 752
rect 878 748 882 752
rect 918 748 922 752
rect 966 748 970 752
rect 1014 748 1018 752
rect 1046 748 1050 752
rect 1062 748 1066 752
rect 102 738 106 742
rect 150 738 154 742
rect 198 738 202 742
rect 390 738 394 742
rect 422 738 426 742
rect 478 738 482 742
rect 510 738 514 742
rect 534 738 538 742
rect 702 738 706 742
rect 726 738 730 742
rect 750 738 754 742
rect 782 738 786 742
rect 838 738 842 742
rect 926 738 930 742
rect 934 738 938 742
rect 958 738 962 742
rect 1006 738 1010 742
rect 1094 747 1098 751
rect 1174 748 1178 752
rect 1206 748 1210 752
rect 1246 748 1250 752
rect 1310 747 1314 751
rect 1382 748 1386 752
rect 1406 748 1410 752
rect 1446 748 1450 752
rect 1078 738 1082 742
rect 1174 738 1178 742
rect 1230 738 1234 742
rect 1278 738 1282 742
rect 1294 738 1298 742
rect 174 728 178 732
rect 190 728 194 732
rect 406 728 410 732
rect 510 728 514 732
rect 710 728 714 732
rect 822 728 826 732
rect 862 728 866 732
rect 118 718 122 722
rect 310 718 314 722
rect 414 718 418 722
rect 742 718 746 722
rect 798 718 802 722
rect 990 718 994 722
rect 1158 718 1162 722
rect 1374 718 1378 722
rect 984 703 988 707
rect 989 703 993 707
rect 994 703 998 707
rect 238 688 242 692
rect 494 688 498 692
rect 534 688 538 692
rect 566 688 570 692
rect 766 688 770 692
rect 902 688 906 692
rect 910 688 914 692
rect 1086 688 1090 692
rect 6 678 10 682
rect 86 678 90 682
rect 614 678 618 682
rect 686 678 690 682
rect 750 678 754 682
rect 798 678 802 682
rect 870 678 874 682
rect 966 678 970 682
rect 1094 678 1098 682
rect 1110 678 1114 682
rect 1134 678 1138 682
rect 1302 678 1306 682
rect 30 668 34 672
rect 182 668 186 672
rect 246 668 250 672
rect 294 668 298 672
rect 374 668 378 672
rect 430 668 434 672
rect 558 668 562 672
rect 590 668 594 672
rect 606 668 610 672
rect 654 668 658 672
rect 662 668 666 672
rect 686 668 690 672
rect 742 668 746 672
rect 766 668 770 672
rect 838 668 842 672
rect 942 668 946 672
rect 1006 668 1010 672
rect 1158 668 1162 672
rect 1238 668 1242 672
rect 1254 668 1258 672
rect 1294 668 1298 672
rect 1358 668 1362 672
rect 1374 668 1378 672
rect 1390 668 1394 672
rect 22 658 26 662
rect 118 659 122 663
rect 182 658 186 662
rect 246 658 250 662
rect 318 658 322 662
rect 350 658 354 662
rect 398 658 402 662
rect 406 658 410 662
rect 454 658 458 662
rect 462 658 466 662
rect 550 658 554 662
rect 582 658 586 662
rect 630 658 634 662
rect 638 658 642 662
rect 670 658 674 662
rect 734 658 738 662
rect 774 658 778 662
rect 886 658 890 662
rect 950 658 954 662
rect 1022 659 1026 663
rect 1150 658 1154 662
rect 1158 658 1162 662
rect 1238 658 1242 662
rect 1270 659 1274 663
rect 1414 658 1418 662
rect 566 648 570 652
rect 710 648 714 652
rect 728 648 732 652
rect 854 648 858 652
rect 918 648 922 652
rect 1182 648 1186 652
rect 822 638 826 642
rect 1150 638 1154 642
rect 422 628 426 632
rect 438 618 442 622
rect 1462 618 1466 622
rect 472 603 476 607
rect 477 603 481 607
rect 482 603 486 607
rect 1414 598 1418 602
rect 278 588 282 592
rect 342 588 346 592
rect 374 588 378 592
rect 478 588 482 592
rect 502 588 506 592
rect 518 588 522 592
rect 1374 588 1378 592
rect 1398 588 1402 592
rect 1422 588 1426 592
rect 1454 588 1458 592
rect 6 578 10 582
rect 1078 578 1082 582
rect 1446 578 1450 582
rect 30 568 34 572
rect 230 568 234 572
rect 270 568 274 572
rect 534 568 538 572
rect 878 568 882 572
rect 894 568 898 572
rect 1150 568 1154 572
rect 102 558 106 562
rect 286 558 290 562
rect 326 558 330 562
rect 614 558 618 562
rect 630 558 634 562
rect 686 558 690 562
rect 702 558 706 562
rect 1006 558 1010 562
rect 1030 558 1034 562
rect 1086 558 1090 562
rect 1166 558 1170 562
rect 1174 558 1178 562
rect 1238 558 1242 562
rect 22 548 26 552
rect 46 548 50 552
rect 70 548 74 552
rect 94 548 98 552
rect 118 548 122 552
rect 166 548 170 552
rect 206 548 210 552
rect 238 548 242 552
rect 270 548 274 552
rect 422 548 426 552
rect 454 548 458 552
rect 470 548 474 552
rect 54 538 58 542
rect 78 538 82 542
rect 94 538 98 542
rect 118 538 122 542
rect 142 538 146 542
rect 158 538 162 542
rect 326 538 330 542
rect 382 538 386 542
rect 414 538 418 542
rect 582 547 586 551
rect 638 548 642 552
rect 654 548 658 552
rect 686 548 690 552
rect 742 548 746 552
rect 838 548 842 552
rect 934 548 938 552
rect 974 548 978 552
rect 1126 548 1130 552
rect 1158 548 1162 552
rect 1174 548 1178 552
rect 1190 548 1194 552
rect 598 538 602 542
rect 646 538 650 542
rect 718 538 722 542
rect 814 538 818 542
rect 854 538 858 542
rect 942 538 946 542
rect 966 538 970 542
rect 1014 538 1018 542
rect 1038 538 1042 542
rect 1062 538 1066 542
rect 1134 538 1138 542
rect 1286 547 1290 551
rect 1382 548 1386 552
rect 1406 548 1410 552
rect 1430 548 1434 552
rect 1470 548 1474 552
rect 1198 538 1202 542
rect 1254 538 1258 542
rect 1294 538 1298 542
rect 54 528 58 532
rect 78 528 82 532
rect 150 528 154 532
rect 190 528 194 532
rect 254 528 258 532
rect 294 528 298 532
rect 350 528 354 532
rect 358 528 362 532
rect 454 528 458 532
rect 510 528 514 532
rect 1054 528 1058 532
rect 1318 528 1322 532
rect 182 518 186 522
rect 390 518 394 522
rect 798 518 802 522
rect 942 518 946 522
rect 1030 518 1034 522
rect 1046 518 1050 522
rect 1094 518 1098 522
rect 1158 518 1162 522
rect 984 503 988 507
rect 989 503 993 507
rect 994 503 998 507
rect 94 488 98 492
rect 166 488 170 492
rect 190 488 194 492
rect 430 488 434 492
rect 470 488 474 492
rect 518 488 522 492
rect 614 488 618 492
rect 1014 488 1018 492
rect 1454 488 1458 492
rect 126 478 130 482
rect 270 478 274 482
rect 334 478 338 482
rect 350 478 354 482
rect 38 468 42 472
rect 118 468 122 472
rect 262 468 266 472
rect 278 468 282 472
rect 326 468 330 472
rect 358 468 362 472
rect 438 478 442 482
rect 494 478 498 482
rect 510 478 514 482
rect 542 478 546 482
rect 774 478 778 482
rect 854 478 858 482
rect 1078 478 1082 482
rect 1110 478 1114 482
rect 1302 478 1306 482
rect 1390 478 1394 482
rect 406 468 410 472
rect 454 468 458 472
rect 462 468 466 472
rect 534 468 538 472
rect 750 468 754 472
rect 822 468 826 472
rect 974 468 978 472
rect 990 468 994 472
rect 1046 468 1050 472
rect 1062 468 1066 472
rect 1078 468 1082 472
rect 1102 468 1106 472
rect 1134 468 1138 472
rect 1142 468 1146 472
rect 1166 468 1170 472
rect 1262 468 1266 472
rect 1270 468 1274 472
rect 1286 468 1290 472
rect 1310 468 1314 472
rect 1358 468 1362 472
rect 46 458 50 462
rect 62 458 66 462
rect 142 458 146 462
rect 190 458 194 462
rect 222 458 226 462
rect 262 458 266 462
rect 318 458 322 462
rect 382 458 386 462
rect 414 458 418 462
rect 558 458 562 462
rect 574 458 578 462
rect 590 458 594 462
rect 598 458 602 462
rect 662 458 666 462
rect 726 458 730 462
rect 758 458 762 462
rect 822 458 826 462
rect 862 458 866 462
rect 1054 458 1058 462
rect 1070 458 1074 462
rect 1126 458 1130 462
rect 1158 458 1162 462
rect 1182 458 1186 462
rect 1222 458 1226 462
rect 1254 458 1258 462
rect 1286 458 1290 462
rect 1342 458 1346 462
rect 1390 459 1394 463
rect 166 448 170 452
rect 198 448 202 452
rect 230 448 234 452
rect 254 448 258 452
rect 430 448 434 452
rect 438 448 442 452
rect 518 448 522 452
rect 942 448 946 452
rect 1086 448 1090 452
rect 1110 448 1114 452
rect 1174 448 1178 452
rect 1230 448 1234 452
rect 1254 448 1258 452
rect 1286 448 1290 452
rect 198 438 202 442
rect 214 438 218 442
rect 382 438 386 442
rect 1190 438 1194 442
rect 1214 438 1218 442
rect 110 418 114 422
rect 294 418 298 422
rect 446 418 450 422
rect 718 418 722 422
rect 918 418 922 422
rect 1182 418 1186 422
rect 472 403 476 407
rect 477 403 481 407
rect 482 403 486 407
rect 230 388 234 392
rect 270 388 274 392
rect 566 388 570 392
rect 814 388 818 392
rect 870 388 874 392
rect 1374 388 1378 392
rect 1398 388 1402 392
rect 1422 388 1426 392
rect 1446 388 1450 392
rect 110 378 114 382
rect 398 378 402 382
rect 654 378 658 382
rect 94 368 98 372
rect 118 368 122 372
rect 390 368 394 372
rect 430 368 434 372
rect 638 368 642 372
rect 1014 368 1018 372
rect 1454 368 1458 372
rect 126 358 130 362
rect 142 358 146 362
rect 182 358 186 362
rect 214 358 218 362
rect 406 358 410 362
rect 590 358 594 362
rect 622 358 626 362
rect 678 358 682 362
rect 710 358 714 362
rect 782 358 786 362
rect 1030 358 1034 362
rect 1126 358 1130 362
rect 1198 358 1202 362
rect 1206 358 1210 362
rect 1238 358 1242 362
rect 1310 358 1314 362
rect 1334 358 1338 362
rect 86 348 90 352
rect 126 348 130 352
rect 190 348 194 352
rect 214 348 218 352
rect 246 348 250 352
rect 262 348 266 352
rect 270 348 274 352
rect 318 348 322 352
rect 374 348 378 352
rect 398 348 402 352
rect 454 348 458 352
rect 462 348 466 352
rect 70 338 74 342
rect 158 338 162 342
rect 166 338 170 342
rect 310 338 314 342
rect 358 338 362 342
rect 502 347 506 351
rect 614 348 618 352
rect 630 348 634 352
rect 654 348 658 352
rect 694 348 698 352
rect 702 348 706 352
rect 726 348 730 352
rect 758 348 762 352
rect 910 348 914 352
rect 950 348 954 352
rect 974 348 978 352
rect 1014 348 1018 352
rect 1038 348 1042 352
rect 1054 348 1058 352
rect 1070 348 1074 352
rect 1086 348 1090 352
rect 1110 348 1114 352
rect 1182 348 1186 352
rect 1222 348 1226 352
rect 1358 348 1362 352
rect 1382 348 1386 352
rect 1406 348 1410 352
rect 1430 348 1434 352
rect 1470 348 1474 352
rect 454 338 458 342
rect 486 338 490 342
rect 574 338 578 342
rect 726 338 730 342
rect 798 338 802 342
rect 846 338 850 342
rect 854 338 858 342
rect 902 338 906 342
rect 998 338 1002 342
rect 1046 338 1050 342
rect 1078 338 1082 342
rect 1102 338 1106 342
rect 1206 338 1210 342
rect 1222 338 1226 342
rect 1254 338 1258 342
rect 1310 338 1314 342
rect 1326 338 1330 342
rect 1350 338 1354 342
rect 54 328 58 332
rect 62 328 66 332
rect 94 328 98 332
rect 238 328 242 332
rect 262 328 266 332
rect 286 328 290 332
rect 302 328 306 332
rect 414 328 418 332
rect 598 328 602 332
rect 630 328 634 332
rect 670 328 674 332
rect 942 328 946 332
rect 1062 328 1066 332
rect 1094 328 1098 332
rect 1158 328 1162 332
rect 1198 328 1202 332
rect 1246 328 1250 332
rect 30 318 34 322
rect 150 318 154 322
rect 174 318 178 322
rect 214 318 218 322
rect 342 318 346 322
rect 582 318 586 322
rect 606 318 610 322
rect 678 318 682 322
rect 750 318 754 322
rect 926 318 930 322
rect 958 318 962 322
rect 1150 318 1154 322
rect 1286 318 1290 322
rect 1310 318 1314 322
rect 1334 318 1338 322
rect 984 303 988 307
rect 989 303 993 307
rect 994 303 998 307
rect 94 288 98 292
rect 302 288 306 292
rect 334 288 338 292
rect 406 288 410 292
rect 518 288 522 292
rect 718 288 722 292
rect 990 288 994 292
rect 1022 288 1026 292
rect 1046 288 1050 292
rect 1230 288 1234 292
rect 1422 288 1426 292
rect 1446 288 1450 292
rect 1454 288 1458 292
rect 198 278 202 282
rect 294 278 298 282
rect 358 278 362 282
rect 446 278 450 282
rect 574 278 578 282
rect 606 278 610 282
rect 750 278 754 282
rect 822 278 826 282
rect 1094 278 1098 282
rect 1134 278 1138 282
rect 1150 278 1154 282
rect 1238 278 1242 282
rect 1278 278 1282 282
rect 1326 278 1330 282
rect 38 268 42 272
rect 190 268 194 272
rect 246 268 250 272
rect 254 268 258 272
rect 270 268 274 272
rect 286 268 290 272
rect 310 268 314 272
rect 326 268 330 272
rect 358 268 362 272
rect 430 268 434 272
rect 486 268 490 272
rect 542 268 546 272
rect 558 268 562 272
rect 606 268 610 272
rect 886 268 890 272
rect 894 268 898 272
rect 942 268 946 272
rect 958 268 962 272
rect 1086 268 1090 272
rect 1102 268 1106 272
rect 1222 268 1226 272
rect 1318 268 1322 272
rect 1374 268 1378 272
rect 38 258 42 262
rect 110 258 114 262
rect 238 258 242 262
rect 246 258 250 262
rect 262 258 266 262
rect 278 258 282 262
rect 374 258 378 262
rect 438 258 442 262
rect 566 258 570 262
rect 598 258 602 262
rect 654 259 658 263
rect 686 258 690 262
rect 758 258 762 262
rect 838 258 842 262
rect 902 258 906 262
rect 950 258 954 262
rect 966 258 970 262
rect 990 258 994 262
rect 1030 258 1034 262
rect 1062 258 1066 262
rect 1094 258 1098 262
rect 1110 258 1114 262
rect 1174 258 1178 262
rect 1182 258 1186 262
rect 1190 258 1194 262
rect 1230 258 1234 262
rect 1366 258 1370 262
rect 1430 258 1434 262
rect 1478 258 1482 262
rect 126 248 130 252
rect 134 248 138 252
rect 174 248 178 252
rect 222 248 226 252
rect 334 248 338 252
rect 398 248 402 252
rect 510 248 514 252
rect 918 248 922 252
rect 982 248 986 252
rect 1054 248 1058 252
rect 214 238 218 242
rect 798 238 802 242
rect 1070 238 1074 242
rect 1126 238 1130 242
rect 1198 238 1202 242
rect 1286 238 1290 242
rect 142 218 146 222
rect 158 218 162 222
rect 238 218 242 222
rect 302 218 306 222
rect 926 218 930 222
rect 1062 218 1066 222
rect 1110 218 1114 222
rect 1190 218 1194 222
rect 472 203 476 207
rect 477 203 481 207
rect 482 203 486 207
rect 22 188 26 192
rect 174 188 178 192
rect 358 188 362 192
rect 430 188 434 192
rect 486 188 490 192
rect 542 188 546 192
rect 614 188 618 192
rect 670 188 674 192
rect 862 188 866 192
rect 878 188 882 192
rect 942 188 946 192
rect 206 178 210 182
rect 974 178 978 182
rect 14 168 18 172
rect 182 168 186 172
rect 270 168 274 172
rect 446 168 450 172
rect 574 168 578 172
rect 606 168 610 172
rect 966 168 970 172
rect 30 158 34 162
rect 102 158 106 162
rect 134 158 138 162
rect 166 158 170 162
rect 222 158 226 162
rect 388 158 392 162
rect 398 158 402 162
rect 438 158 442 162
rect 446 158 450 162
rect 494 158 498 162
rect 590 158 594 162
rect 678 158 682 162
rect 886 158 890 162
rect 1006 158 1010 162
rect 1070 158 1074 162
rect 1238 158 1242 162
rect 22 148 26 152
rect 62 148 66 152
rect 150 148 154 152
rect 174 148 178 152
rect 206 148 210 152
rect 238 148 242 152
rect 262 148 266 152
rect 270 148 274 152
rect 286 148 290 152
rect 294 148 298 152
rect 350 148 354 152
rect 374 148 378 152
rect 382 148 386 152
rect 398 148 402 152
rect 414 148 418 152
rect 454 148 458 152
rect 494 148 498 152
rect 526 148 530 152
rect 542 148 546 152
rect 558 148 562 152
rect 566 148 570 152
rect 598 148 602 152
rect 630 148 634 152
rect 718 148 722 152
rect 806 148 810 152
rect 918 148 922 152
rect 974 148 978 152
rect 998 148 1002 152
rect 1022 148 1026 152
rect 1078 148 1082 152
rect 1086 148 1090 152
rect 1126 148 1130 152
rect 1134 148 1138 152
rect 1158 148 1162 152
rect 1166 148 1170 152
rect 1206 148 1210 152
rect 1342 148 1346 152
rect 1390 147 1394 151
rect 38 138 42 142
rect 86 138 90 142
rect 126 138 130 142
rect 158 138 162 142
rect 198 138 202 142
rect 230 138 234 142
rect 262 138 266 142
rect 302 138 306 142
rect 374 138 378 142
rect 422 138 426 142
rect 510 138 514 142
rect 518 138 522 142
rect 550 138 554 142
rect 574 138 578 142
rect 638 138 642 142
rect 702 138 706 142
rect 726 138 730 142
rect 798 138 802 142
rect 870 138 874 142
rect 910 138 914 142
rect 1030 138 1034 142
rect 1078 138 1082 142
rect 1126 138 1130 142
rect 1182 138 1186 142
rect 1214 138 1218 142
rect 1222 138 1226 142
rect 1246 138 1250 142
rect 1254 138 1258 142
rect 1302 138 1306 142
rect 1310 138 1314 142
rect 1358 138 1362 142
rect 1374 138 1378 142
rect 1438 138 1442 142
rect 46 128 50 132
rect 238 128 242 132
rect 286 128 290 132
rect 318 128 322 132
rect 342 128 346 132
rect 414 128 418 132
rect 638 128 642 132
rect 694 128 698 132
rect 718 128 722 132
rect 734 128 738 132
rect 902 128 906 132
rect 1038 128 1042 132
rect 1102 128 1106 132
rect 1110 128 1114 132
rect 1198 128 1202 132
rect 1230 128 1234 132
rect 1390 128 1394 132
rect 54 118 58 122
rect 334 118 338 122
rect 862 118 866 122
rect 878 118 882 122
rect 1126 118 1130 122
rect 1190 118 1194 122
rect 1286 118 1290 122
rect 1470 118 1474 122
rect 984 103 988 107
rect 989 103 993 107
rect 994 103 998 107
rect 46 88 50 92
rect 134 88 138 92
rect 190 88 194 92
rect 254 88 258 92
rect 318 88 322 92
rect 502 88 506 92
rect 574 88 578 92
rect 590 88 594 92
rect 718 88 722 92
rect 870 88 874 92
rect 894 88 898 92
rect 918 88 922 92
rect 1070 88 1074 92
rect 1110 88 1114 92
rect 1326 88 1330 92
rect 1422 88 1426 92
rect 1446 88 1450 92
rect 1454 88 1458 92
rect 62 78 66 82
rect 70 78 74 82
rect 118 78 122 82
rect 142 78 146 82
rect 198 78 202 82
rect 238 78 242 82
rect 294 78 298 82
rect 326 78 330 82
rect 382 78 386 82
rect 398 78 402 82
rect 470 78 474 82
rect 486 78 490 82
rect 550 78 554 82
rect 582 78 586 82
rect 838 78 842 82
rect 854 78 858 82
rect 886 78 890 82
rect 46 68 50 72
rect 94 68 98 72
rect 190 68 194 72
rect 222 68 226 72
rect 230 68 234 72
rect 318 68 322 72
rect 358 68 362 72
rect 390 68 394 72
rect 510 68 514 72
rect 670 68 674 72
rect 686 68 690 72
rect 734 68 738 72
rect 742 68 746 72
rect 806 68 810 72
rect 814 68 818 72
rect 830 68 834 72
rect 878 68 882 72
rect 910 68 914 72
rect 1006 78 1010 82
rect 1062 78 1066 82
rect 1118 78 1122 82
rect 1142 78 1146 82
rect 934 68 938 72
rect 982 66 986 70
rect 1014 68 1018 72
rect 1062 68 1066 72
rect 1102 68 1106 72
rect 1230 68 1234 72
rect 1246 68 1250 72
rect 1342 68 1346 72
rect 1390 68 1394 72
rect 94 58 98 62
rect 198 58 202 62
rect 270 58 274 62
rect 278 58 282 62
rect 310 58 314 62
rect 366 58 370 62
rect 414 58 418 62
rect 446 58 450 62
rect 454 58 458 62
rect 470 58 474 62
rect 526 58 530 62
rect 534 58 538 62
rect 558 58 562 62
rect 654 59 658 63
rect 854 58 858 62
rect 918 58 922 62
rect 942 58 946 62
rect 1054 58 1058 62
rect 1126 58 1130 62
rect 1158 58 1162 62
rect 1230 58 1234 62
rect 1262 59 1266 63
rect 1358 59 1362 63
rect 1430 58 1434 62
rect 1470 58 1474 62
rect 214 48 218 52
rect 246 48 250 52
rect 254 48 258 52
rect 750 48 754 52
rect 814 48 818 52
rect 862 48 866 52
rect 1078 48 1082 52
rect 1174 48 1178 52
rect 294 38 298 42
rect 774 38 778 42
rect 942 38 946 42
rect 472 3 476 7
rect 477 3 481 7
rect 482 3 486 7
<< metal2 >>
rect 158 1192 161 1208
rect 230 1192 233 1198
rect 310 1192 313 1198
rect 334 1192 337 1208
rect 186 1188 190 1191
rect 210 1178 214 1181
rect 42 1148 46 1151
rect 102 1132 105 1168
rect 238 1152 241 1168
rect 350 1162 353 1231
rect 366 1202 369 1231
rect 382 1228 393 1231
rect 406 1228 417 1231
rect 382 1192 385 1228
rect 390 1192 393 1198
rect 414 1192 417 1228
rect 422 1228 433 1231
rect 422 1192 425 1228
rect 434 1188 438 1191
rect 446 1181 449 1231
rect 454 1228 473 1231
rect 478 1228 489 1231
rect 454 1192 457 1228
rect 478 1221 481 1228
rect 462 1218 481 1221
rect 462 1202 465 1218
rect 476 1203 477 1207
rect 481 1203 482 1207
rect 486 1203 488 1207
rect 494 1191 497 1208
rect 482 1188 497 1191
rect 438 1178 449 1181
rect 526 1182 529 1231
rect 542 1202 545 1231
rect 566 1202 569 1231
rect 582 1202 585 1231
rect 606 1212 609 1231
rect 622 1211 625 1231
rect 646 1212 649 1231
rect 622 1208 633 1211
rect 366 1152 369 1158
rect 118 1142 121 1148
rect 106 1128 110 1131
rect 30 1082 33 1128
rect 94 1082 97 1088
rect 106 1078 110 1081
rect 134 1072 137 1148
rect 118 1062 121 1068
rect 134 1062 137 1068
rect 50 1058 54 1061
rect 62 952 65 1058
rect 98 988 102 991
rect 58 948 62 951
rect 38 942 41 948
rect 118 942 121 948
rect 30 882 33 928
rect 98 888 102 891
rect 118 862 121 868
rect 134 862 137 938
rect 142 892 145 1148
rect 166 1082 169 1148
rect 190 1132 193 1148
rect 206 1082 209 1148
rect 214 1092 217 1148
rect 238 1072 241 1138
rect 174 1062 177 1068
rect 166 962 169 1058
rect 182 972 185 1018
rect 166 952 169 958
rect 198 951 201 968
rect 222 952 225 1068
rect 254 1062 257 1118
rect 262 992 265 1148
rect 270 1142 273 1148
rect 286 1142 289 1148
rect 318 1132 321 1148
rect 290 1128 294 1131
rect 270 1062 273 1068
rect 286 992 289 1118
rect 302 1092 305 1128
rect 350 1072 353 1118
rect 350 1062 353 1068
rect 358 1062 361 1068
rect 326 952 329 968
rect 350 952 353 1058
rect 42 858 46 861
rect 62 752 65 758
rect 94 752 97 768
rect 150 752 153 918
rect 230 882 233 888
rect 270 882 273 948
rect 242 878 246 881
rect 198 862 201 868
rect 254 862 257 868
rect 278 862 281 948
rect 310 882 313 888
rect 294 862 297 868
rect 310 862 313 868
rect 178 858 182 861
rect 198 762 201 858
rect 342 852 345 859
rect 366 852 369 1148
rect 374 1102 377 1148
rect 398 1112 401 1148
rect 382 992 385 1108
rect 422 1092 425 1148
rect 438 1122 441 1178
rect 630 1172 633 1208
rect 662 1182 665 1231
rect 686 1192 689 1231
rect 694 1192 697 1208
rect 686 1172 689 1178
rect 734 1172 737 1178
rect 666 1168 670 1171
rect 506 1158 510 1161
rect 622 1152 625 1168
rect 634 1158 638 1161
rect 402 1088 406 1091
rect 422 1082 425 1088
rect 426 1058 430 1061
rect 394 968 398 971
rect 406 952 409 1058
rect 446 972 449 1148
rect 482 1138 486 1141
rect 514 1138 518 1141
rect 502 1081 505 1118
rect 550 1092 553 1147
rect 502 1078 510 1081
rect 482 1068 486 1071
rect 538 1068 542 1071
rect 566 1062 569 1068
rect 454 982 457 1058
rect 526 1052 529 1058
rect 534 1032 537 1058
rect 394 948 398 951
rect 386 928 390 931
rect 414 892 417 968
rect 422 932 425 938
rect 430 932 433 968
rect 450 948 454 951
rect 442 928 446 931
rect 402 888 406 891
rect 38 732 41 748
rect 6 682 9 688
rect 22 662 25 668
rect 30 662 33 668
rect 6 582 9 588
rect 30 562 33 568
rect 26 548 30 551
rect 46 542 49 548
rect 54 542 57 548
rect 54 522 57 528
rect 22 192 25 218
rect 30 201 33 318
rect 38 272 41 468
rect 62 462 65 748
rect 150 742 153 748
rect 102 722 105 738
rect 174 732 177 748
rect 86 682 89 718
rect 118 663 121 718
rect 182 672 185 758
rect 206 752 209 818
rect 230 792 233 838
rect 218 748 222 751
rect 194 738 198 741
rect 190 722 193 728
rect 262 712 265 748
rect 286 712 289 748
rect 314 718 318 721
rect 238 672 241 688
rect 294 672 297 678
rect 242 668 246 671
rect 318 662 321 708
rect 118 658 121 659
rect 186 658 190 661
rect 242 658 246 661
rect 322 658 326 661
rect 342 592 345 828
rect 374 812 377 858
rect 374 751 377 768
rect 422 752 425 778
rect 374 662 377 668
rect 354 658 358 661
rect 374 592 377 648
rect 282 588 286 591
rect 230 572 233 578
rect 254 562 257 578
rect 266 568 270 571
rect 70 552 73 558
rect 102 552 105 558
rect 118 552 121 558
rect 206 552 209 558
rect 90 548 94 551
rect 170 548 174 551
rect 74 538 78 541
rect 94 532 97 538
rect 118 532 121 538
rect 82 528 86 531
rect 98 488 102 491
rect 126 482 129 528
rect 118 472 121 478
rect 38 222 41 258
rect 46 232 49 458
rect 110 402 113 418
rect 54 332 57 398
rect 110 382 113 388
rect 98 368 102 371
rect 114 368 118 371
rect 126 362 129 478
rect 142 472 145 538
rect 158 532 161 538
rect 150 492 153 528
rect 166 492 169 518
rect 142 462 145 468
rect 142 362 145 368
rect 150 352 153 488
rect 166 442 169 448
rect 130 348 134 351
rect 86 342 89 348
rect 30 198 41 201
rect 14 162 17 168
rect 30 162 33 188
rect 26 148 30 151
rect 38 142 41 198
rect 62 162 65 328
rect 70 322 73 338
rect 86 161 89 338
rect 98 328 102 331
rect 94 292 97 328
rect 110 262 113 348
rect 158 342 161 358
rect 174 351 177 548
rect 182 462 185 518
rect 190 502 193 528
rect 190 492 193 498
rect 190 462 193 468
rect 198 452 201 478
rect 230 472 233 538
rect 238 522 241 548
rect 254 532 257 558
rect 270 522 273 548
rect 254 471 257 498
rect 266 478 270 481
rect 278 472 281 528
rect 254 468 262 471
rect 166 348 177 351
rect 182 362 185 448
rect 214 442 217 458
rect 222 452 225 458
rect 230 452 233 468
rect 254 442 257 448
rect 166 342 169 348
rect 134 252 137 268
rect 126 242 129 248
rect 142 192 145 218
rect 86 158 97 161
rect 106 158 110 161
rect 46 92 49 128
rect 54 122 57 158
rect 62 132 65 148
rect 70 82 73 158
rect 86 142 89 148
rect 50 68 54 71
rect 62 62 65 78
rect 70 -22 73 78
rect 94 72 97 158
rect 118 82 121 168
rect 134 162 137 168
rect 126 122 129 138
rect 134 92 137 148
rect 142 82 145 178
rect 150 152 153 318
rect 158 272 161 338
rect 166 332 169 338
rect 182 332 185 358
rect 190 352 193 398
rect 166 292 169 328
rect 178 318 182 321
rect 198 282 201 438
rect 230 392 233 428
rect 214 362 217 378
rect 214 352 217 358
rect 262 352 265 458
rect 270 392 273 458
rect 286 442 289 558
rect 294 492 297 528
rect 294 372 297 418
rect 250 348 254 351
rect 246 342 249 348
rect 242 328 246 331
rect 186 268 190 271
rect 198 252 201 278
rect 170 248 174 251
rect 158 182 161 218
rect 174 192 177 228
rect 206 191 209 298
rect 214 272 217 318
rect 222 282 225 328
rect 222 252 225 278
rect 246 272 249 288
rect 262 282 265 328
rect 254 272 257 278
rect 270 272 273 348
rect 302 342 305 578
rect 390 572 393 738
rect 422 732 425 738
rect 410 728 414 731
rect 398 662 401 668
rect 406 592 409 658
rect 414 582 417 718
rect 430 672 433 808
rect 438 742 441 768
rect 462 762 465 1018
rect 476 1003 477 1007
rect 481 1003 482 1007
rect 486 1003 488 1007
rect 526 962 529 1018
rect 574 1002 577 1148
rect 622 1142 625 1148
rect 638 1142 641 1148
rect 582 1082 585 1128
rect 618 1118 622 1121
rect 594 1058 598 1061
rect 582 992 585 1058
rect 606 992 609 1078
rect 614 1062 617 1108
rect 626 1068 630 1071
rect 614 1052 617 1058
rect 630 1022 633 1058
rect 586 968 590 971
rect 478 952 481 958
rect 534 952 537 958
rect 566 952 569 968
rect 522 948 526 951
rect 522 938 526 941
rect 554 938 558 941
rect 498 928 502 931
rect 478 863 481 868
rect 510 862 513 918
rect 566 872 569 878
rect 530 868 534 871
rect 590 862 593 878
rect 478 858 481 859
rect 550 852 553 858
rect 606 832 609 988
rect 638 942 641 998
rect 638 872 641 938
rect 646 892 649 1148
rect 670 1122 673 1148
rect 710 1102 713 1148
rect 718 1142 721 1158
rect 742 1142 745 1158
rect 750 1152 753 1208
rect 790 1172 793 1178
rect 758 1152 761 1168
rect 774 1162 777 1168
rect 798 1161 801 1198
rect 862 1182 865 1231
rect 790 1158 801 1161
rect 766 1152 769 1158
rect 750 1112 753 1138
rect 686 1092 689 1098
rect 766 1072 769 1138
rect 782 1131 785 1148
rect 790 1142 793 1158
rect 862 1151 865 1158
rect 814 1142 817 1148
rect 782 1128 793 1131
rect 790 1092 793 1128
rect 662 1062 665 1068
rect 782 1062 785 1078
rect 798 1062 801 1088
rect 806 1082 809 1138
rect 806 1062 809 1078
rect 822 1072 825 1148
rect 886 1142 889 1231
rect 902 1192 905 1231
rect 830 1122 833 1138
rect 846 1132 849 1138
rect 926 1132 929 1231
rect 942 1172 945 1231
rect 966 1182 969 1231
rect 982 1192 985 1231
rect 1022 1202 1025 1231
rect 1038 1212 1041 1231
rect 938 1148 942 1151
rect 942 1132 945 1138
rect 950 1132 953 1178
rect 982 1152 985 1158
rect 1038 1152 1041 1158
rect 1034 1148 1038 1151
rect 926 1112 929 1118
rect 830 1062 833 1068
rect 654 1042 657 1048
rect 718 1002 721 1058
rect 742 1052 745 1058
rect 830 1052 833 1058
rect 838 1052 841 1078
rect 862 1072 865 1098
rect 894 1092 897 1098
rect 902 1081 905 1098
rect 894 1078 905 1081
rect 910 1082 913 1088
rect 854 1062 857 1068
rect 846 1048 848 1051
rect 790 1012 793 1018
rect 654 932 657 947
rect 670 862 673 938
rect 686 932 689 968
rect 718 962 721 998
rect 766 962 769 998
rect 782 952 785 988
rect 806 961 809 1018
rect 830 992 833 1048
rect 846 972 849 1048
rect 802 958 809 961
rect 830 962 833 968
rect 738 948 742 951
rect 826 948 830 951
rect 702 942 705 948
rect 722 938 726 941
rect 738 938 742 941
rect 686 882 689 888
rect 702 872 705 938
rect 722 928 726 931
rect 750 912 753 948
rect 718 892 721 898
rect 782 892 785 938
rect 790 892 793 948
rect 802 938 806 941
rect 798 922 801 928
rect 814 922 817 948
rect 846 942 849 958
rect 862 942 865 947
rect 710 872 713 878
rect 726 862 729 868
rect 734 862 737 878
rect 798 872 801 878
rect 476 803 477 807
rect 481 803 482 807
rect 486 803 488 807
rect 486 752 489 778
rect 494 758 502 761
rect 450 748 454 751
rect 478 732 481 738
rect 494 692 497 758
rect 510 752 513 808
rect 614 792 617 858
rect 622 802 625 818
rect 546 768 550 771
rect 610 768 614 771
rect 558 762 561 768
rect 570 758 574 761
rect 514 738 518 741
rect 422 632 425 638
rect 322 558 326 561
rect 330 538 334 541
rect 358 532 361 558
rect 382 542 385 548
rect 422 542 425 548
rect 350 522 353 528
rect 318 452 321 458
rect 326 432 329 468
rect 334 452 337 478
rect 310 342 313 398
rect 302 332 305 338
rect 238 262 241 268
rect 278 262 281 308
rect 286 302 289 328
rect 294 321 297 328
rect 294 318 305 321
rect 302 292 305 318
rect 298 278 302 281
rect 234 258 238 261
rect 266 258 270 261
rect 214 242 217 248
rect 198 188 209 191
rect 238 192 241 218
rect 166 152 169 158
rect 174 152 177 178
rect 150 112 153 148
rect 162 138 166 141
rect 182 102 185 168
rect 198 142 201 188
rect 210 178 214 181
rect 222 152 225 158
rect 210 148 214 151
rect 198 122 201 138
rect 194 88 198 91
rect 202 78 206 81
rect 190 72 193 78
rect 222 72 225 148
rect 230 142 233 168
rect 238 152 241 168
rect 246 142 249 258
rect 278 242 281 258
rect 238 122 241 128
rect 254 92 257 238
rect 286 192 289 268
rect 294 182 297 278
rect 310 272 313 328
rect 318 322 321 348
rect 334 292 337 438
rect 350 402 353 478
rect 358 472 361 478
rect 382 472 385 538
rect 414 532 417 538
rect 394 518 398 521
rect 430 492 433 658
rect 454 652 457 658
rect 438 502 441 618
rect 454 542 457 548
rect 462 542 465 658
rect 476 603 477 607
rect 481 603 482 607
rect 486 603 488 607
rect 502 592 505 708
rect 510 702 513 728
rect 526 722 529 748
rect 518 592 521 698
rect 534 692 537 738
rect 542 732 545 748
rect 574 742 577 748
rect 582 742 585 768
rect 622 762 625 798
rect 646 792 649 818
rect 634 768 638 771
rect 742 762 745 798
rect 650 758 654 761
rect 594 748 598 751
rect 614 742 617 748
rect 646 742 649 748
rect 670 742 673 748
rect 566 692 569 728
rect 606 672 609 718
rect 614 702 617 708
rect 614 682 617 698
rect 562 668 566 671
rect 594 668 598 671
rect 606 662 609 668
rect 554 658 558 661
rect 586 658 590 661
rect 566 592 569 648
rect 614 602 617 678
rect 630 662 633 678
rect 638 662 641 738
rect 686 682 689 758
rect 702 742 705 758
rect 726 742 729 748
rect 750 742 753 868
rect 814 862 817 888
rect 766 812 769 858
rect 786 848 790 851
rect 814 842 817 848
rect 822 842 825 928
rect 846 892 849 918
rect 770 768 774 771
rect 758 761 761 768
rect 758 758 769 761
rect 714 728 718 731
rect 726 702 729 738
rect 662 672 665 678
rect 686 672 689 678
rect 742 672 745 718
rect 750 712 753 738
rect 750 682 753 708
rect 758 702 761 748
rect 766 692 769 758
rect 782 742 785 838
rect 814 782 817 818
rect 838 812 841 878
rect 870 862 873 1068
rect 878 1062 881 1068
rect 878 912 881 1058
rect 894 1052 897 1078
rect 902 1052 905 1068
rect 918 1052 921 1058
rect 942 1042 945 1058
rect 930 1038 934 1041
rect 950 1022 953 1068
rect 958 1042 961 1058
rect 966 1052 969 1148
rect 988 1103 989 1107
rect 993 1103 994 1107
rect 998 1103 1000 1107
rect 1006 1071 1009 1138
rect 998 1068 1009 1071
rect 926 992 929 1008
rect 958 962 961 968
rect 966 952 969 1048
rect 998 962 1001 1068
rect 1014 1062 1017 1128
rect 1022 1062 1025 1098
rect 1038 1082 1041 1088
rect 1030 1062 1033 1068
rect 1038 1062 1041 1078
rect 1046 1062 1049 1178
rect 1062 1172 1065 1231
rect 1078 1228 1089 1231
rect 1078 1172 1081 1208
rect 1054 1132 1057 1168
rect 1086 1152 1089 1228
rect 1102 1192 1105 1231
rect 1118 1212 1121 1231
rect 1110 1172 1113 1198
rect 1142 1182 1145 1231
rect 1158 1228 1169 1231
rect 1150 1172 1153 1188
rect 1166 1182 1169 1228
rect 1182 1202 1185 1231
rect 1198 1212 1201 1231
rect 1222 1182 1225 1231
rect 1238 1202 1241 1231
rect 1206 1172 1209 1178
rect 1222 1162 1225 1168
rect 1126 1152 1129 1158
rect 1174 1152 1177 1158
rect 1134 1142 1137 1148
rect 1106 1138 1110 1141
rect 1130 1138 1134 1141
rect 1054 1092 1057 1098
rect 1062 1072 1065 1138
rect 1070 1082 1073 1118
rect 1078 1072 1081 1138
rect 1158 1132 1161 1138
rect 1098 1118 1102 1121
rect 1118 1091 1121 1118
rect 1142 1112 1145 1118
rect 1110 1088 1121 1091
rect 1078 1062 1081 1068
rect 1006 1052 1009 1058
rect 1070 1052 1073 1058
rect 1086 1042 1089 1068
rect 1094 1052 1097 1058
rect 1110 1052 1113 1088
rect 1118 1072 1121 1078
rect 1134 1062 1137 1088
rect 1142 1062 1145 1098
rect 1166 1062 1169 1068
rect 1174 1062 1177 1148
rect 1222 1142 1225 1148
rect 1246 1142 1249 1148
rect 1262 1142 1265 1231
rect 1278 1212 1281 1231
rect 1302 1228 1313 1231
rect 1270 1172 1273 1188
rect 1194 1128 1198 1131
rect 1190 1071 1193 1118
rect 1214 1092 1217 1118
rect 1182 1068 1193 1071
rect 1206 1072 1209 1078
rect 1182 1052 1185 1068
rect 1194 1058 1198 1061
rect 886 862 889 888
rect 862 832 865 858
rect 870 852 873 858
rect 810 768 814 771
rect 802 758 806 761
rect 822 752 825 798
rect 830 752 833 758
rect 838 752 841 808
rect 870 762 873 798
rect 894 792 897 868
rect 910 862 913 948
rect 922 918 926 921
rect 918 882 921 918
rect 934 902 937 938
rect 942 912 945 948
rect 994 918 998 921
rect 930 878 934 881
rect 946 858 950 861
rect 910 812 913 858
rect 958 852 961 918
rect 988 903 989 907
rect 993 903 994 907
rect 998 903 1000 907
rect 974 882 977 888
rect 966 862 969 868
rect 982 862 985 868
rect 966 852 969 858
rect 918 848 926 851
rect 942 848 950 851
rect 918 822 921 848
rect 930 828 934 831
rect 942 792 945 848
rect 902 772 905 778
rect 890 768 894 771
rect 854 758 862 761
rect 834 738 838 741
rect 782 732 785 738
rect 822 732 825 738
rect 798 682 801 718
rect 846 692 849 748
rect 854 732 857 758
rect 878 752 881 768
rect 922 748 926 751
rect 862 732 865 738
rect 750 672 753 678
rect 650 668 654 671
rect 834 668 838 671
rect 734 662 737 668
rect 638 652 641 658
rect 670 642 673 658
rect 766 652 769 668
rect 778 658 782 661
rect 854 652 857 698
rect 902 692 905 718
rect 910 682 913 688
rect 866 678 870 681
rect 706 648 710 651
rect 726 648 728 651
rect 482 588 486 591
rect 530 568 534 571
rect 614 562 617 588
rect 582 551 585 558
rect 630 552 633 558
rect 638 552 641 598
rect 450 528 454 531
rect 442 478 446 481
rect 454 472 457 528
rect 470 492 473 548
rect 646 542 649 588
rect 654 552 657 598
rect 726 592 729 648
rect 826 638 830 641
rect 686 562 689 568
rect 702 562 705 568
rect 682 548 686 551
rect 718 542 721 548
rect 514 528 521 531
rect 518 492 521 528
rect 462 472 465 488
rect 542 482 545 488
rect 498 478 502 481
rect 510 472 513 478
rect 378 458 382 461
rect 382 442 385 448
rect 386 368 390 371
rect 398 362 401 378
rect 406 372 409 468
rect 414 452 417 458
rect 438 452 441 468
rect 454 452 457 468
rect 514 448 518 451
rect 430 372 433 448
rect 534 442 537 468
rect 558 452 561 458
rect 446 422 449 428
rect 476 403 477 407
rect 481 403 482 407
rect 486 403 488 407
rect 374 342 377 348
rect 354 338 358 341
rect 346 318 350 321
rect 322 268 326 271
rect 310 262 313 268
rect 330 248 334 251
rect 270 161 273 168
rect 262 158 273 161
rect 262 152 265 158
rect 270 142 273 148
rect 262 132 265 138
rect 242 78 246 81
rect 198 62 201 68
rect 94 52 97 58
rect 214 52 217 58
rect 230 -22 233 68
rect 278 62 281 178
rect 294 152 297 158
rect 286 132 289 148
rect 294 82 297 148
rect 302 142 305 218
rect 342 182 345 318
rect 398 282 401 348
rect 406 292 409 358
rect 414 322 417 328
rect 358 272 361 278
rect 358 192 361 268
rect 374 262 377 278
rect 422 272 425 368
rect 454 352 457 378
rect 502 351 505 358
rect 450 338 454 341
rect 426 268 430 271
rect 446 262 449 278
rect 378 258 382 261
rect 430 258 438 261
rect 394 248 398 251
rect 318 132 321 138
rect 326 102 329 178
rect 342 132 345 168
rect 350 152 353 188
rect 390 162 393 168
rect 392 158 393 162
rect 398 162 401 248
rect 430 192 433 258
rect 446 182 449 258
rect 446 172 449 178
rect 454 162 457 338
rect 402 148 406 151
rect 374 142 377 148
rect 382 132 385 148
rect 414 132 417 148
rect 422 142 425 158
rect 438 142 441 158
rect 446 152 449 158
rect 454 142 457 148
rect 462 142 465 348
rect 486 342 489 348
rect 522 288 526 291
rect 558 272 561 438
rect 566 392 569 538
rect 598 532 601 538
rect 614 492 617 538
rect 574 462 577 478
rect 590 462 593 468
rect 602 458 606 461
rect 722 458 726 461
rect 662 442 665 458
rect 570 388 574 391
rect 658 378 662 381
rect 590 362 593 378
rect 638 372 641 378
rect 630 362 633 368
rect 574 342 577 358
rect 614 342 617 348
rect 574 332 577 338
rect 570 278 574 281
rect 490 268 497 271
rect 538 268 542 271
rect 476 203 477 207
rect 481 203 482 207
rect 486 203 488 207
rect 494 191 497 268
rect 558 262 561 268
rect 510 242 513 248
rect 490 188 497 191
rect 542 192 545 248
rect 566 242 569 258
rect 318 92 321 98
rect 310 62 313 88
rect 326 82 329 98
rect 334 92 337 118
rect 378 78 382 81
rect 390 72 393 98
rect 398 82 401 88
rect 322 68 326 71
rect 354 68 358 71
rect 462 71 465 138
rect 470 82 473 158
rect 486 82 489 178
rect 494 162 497 168
rect 498 148 502 151
rect 510 142 513 178
rect 566 152 569 238
rect 582 192 585 318
rect 598 312 601 328
rect 606 282 609 318
rect 610 268 614 271
rect 598 252 601 258
rect 614 192 617 248
rect 622 182 625 358
rect 630 352 633 358
rect 650 348 654 351
rect 670 342 673 448
rect 678 362 681 418
rect 718 412 721 418
rect 710 362 713 368
rect 694 352 697 358
rect 726 352 729 458
rect 742 452 745 548
rect 750 472 753 618
rect 878 572 881 668
rect 886 662 889 678
rect 918 662 921 748
rect 926 732 929 738
rect 934 702 937 738
rect 942 672 945 738
rect 950 722 953 838
rect 982 762 985 818
rect 1014 761 1017 1018
rect 1030 992 1033 1018
rect 1126 982 1129 1018
rect 1142 962 1145 968
rect 1046 952 1049 958
rect 1062 952 1065 958
rect 1158 952 1161 1018
rect 1022 932 1025 948
rect 1046 922 1049 948
rect 1054 942 1057 948
rect 1086 942 1089 948
rect 1078 932 1081 938
rect 1086 922 1089 928
rect 1030 892 1033 918
rect 1022 862 1025 868
rect 1046 862 1049 898
rect 1054 872 1057 918
rect 1102 902 1105 948
rect 1110 942 1113 948
rect 1158 932 1161 938
rect 1166 932 1169 988
rect 1182 942 1185 978
rect 1190 952 1193 1058
rect 1198 972 1201 1018
rect 1206 952 1209 1058
rect 1214 1052 1217 1068
rect 1222 1062 1225 1138
rect 1230 1062 1233 1068
rect 1238 1052 1241 1118
rect 1246 1062 1249 1068
rect 1254 1062 1257 1138
rect 1262 1072 1265 1078
rect 1270 1052 1273 1118
rect 1286 1081 1289 1198
rect 1294 1092 1297 1148
rect 1310 1092 1313 1228
rect 1318 1212 1321 1231
rect 1342 1202 1345 1231
rect 1322 1188 1326 1191
rect 1350 1191 1353 1208
rect 1346 1188 1353 1191
rect 1322 1148 1326 1151
rect 1346 1148 1350 1151
rect 1286 1078 1297 1081
rect 1278 1052 1281 1058
rect 1214 1032 1217 1048
rect 1230 992 1233 1048
rect 1294 992 1297 1078
rect 1318 992 1321 1138
rect 1326 1062 1329 1148
rect 1358 1142 1361 1231
rect 1366 1192 1369 1208
rect 1366 1081 1369 1178
rect 1382 1162 1385 1231
rect 1398 1212 1401 1231
rect 1414 1228 1425 1231
rect 1430 1228 1441 1231
rect 1414 1192 1417 1228
rect 1430 1202 1433 1228
rect 1438 1192 1441 1208
rect 1462 1192 1465 1231
rect 1478 1212 1481 1231
rect 1390 1182 1393 1188
rect 1378 1148 1382 1151
rect 1418 1148 1422 1151
rect 1374 1092 1377 1128
rect 1398 1092 1401 1148
rect 1414 1092 1417 1138
rect 1366 1078 1377 1081
rect 1358 1062 1361 1068
rect 1350 1051 1353 1058
rect 1350 1048 1361 1051
rect 1222 962 1225 968
rect 1246 952 1249 988
rect 1278 952 1281 958
rect 1342 952 1345 1048
rect 1358 992 1361 1048
rect 1374 992 1377 1078
rect 1382 1052 1385 1058
rect 1398 992 1401 1078
rect 1430 1062 1433 1148
rect 1438 1092 1441 1168
rect 1446 1071 1449 1148
rect 1478 1092 1481 1158
rect 1438 1068 1449 1071
rect 1438 1012 1441 1068
rect 1486 1062 1489 1118
rect 1450 1058 1454 1061
rect 1358 962 1361 988
rect 1438 952 1441 958
rect 1462 952 1465 958
rect 1258 948 1262 951
rect 1314 948 1318 951
rect 1330 948 1334 951
rect 1410 948 1414 951
rect 1062 872 1065 878
rect 1094 872 1097 878
rect 1146 868 1150 871
rect 1030 802 1033 818
rect 1046 812 1049 858
rect 1054 842 1057 868
rect 1086 862 1089 868
rect 1134 862 1137 868
rect 1070 852 1073 858
rect 1102 852 1105 858
rect 1158 852 1161 868
rect 1086 842 1089 848
rect 1086 822 1089 838
rect 1046 762 1049 808
rect 1166 792 1169 908
rect 1174 872 1177 918
rect 1190 892 1193 948
rect 1198 902 1201 938
rect 1238 922 1241 928
rect 1182 872 1185 878
rect 1178 858 1182 861
rect 1198 792 1201 878
rect 1222 872 1225 918
rect 1218 859 1222 861
rect 1214 858 1222 859
rect 1238 822 1241 918
rect 1246 862 1249 868
rect 1270 862 1273 918
rect 1278 842 1281 848
rect 1282 838 1286 841
rect 1062 762 1065 768
rect 1014 758 1025 761
rect 966 742 969 748
rect 1014 742 1017 748
rect 958 732 961 738
rect 1006 732 1009 738
rect 994 718 998 721
rect 1014 712 1017 738
rect 988 703 989 707
rect 993 703 994 707
rect 998 703 1000 707
rect 966 682 969 688
rect 918 652 921 658
rect 942 652 945 668
rect 1006 662 1009 668
rect 1022 663 1025 758
rect 1206 752 1209 808
rect 1222 762 1225 768
rect 1046 722 1049 748
rect 1062 742 1065 748
rect 1178 748 1182 751
rect 1250 748 1254 751
rect 1094 742 1097 747
rect 1294 742 1297 868
rect 1310 863 1313 868
rect 1342 862 1345 948
rect 1390 892 1393 948
rect 1430 862 1433 948
rect 1310 858 1313 859
rect 1402 858 1406 861
rect 1342 792 1345 858
rect 1378 818 1382 821
rect 1398 792 1401 798
rect 1406 752 1409 818
rect 1422 782 1425 788
rect 1438 751 1441 948
rect 1462 892 1465 918
rect 1478 842 1481 858
rect 1486 812 1489 898
rect 1438 748 1446 751
rect 1310 742 1313 747
rect 1226 738 1230 741
rect 1078 672 1081 738
rect 1158 712 1161 718
rect 1174 712 1177 738
rect 1086 692 1089 698
rect 1090 678 1094 681
rect 1110 672 1113 678
rect 1022 658 1025 659
rect 950 592 953 658
rect 1134 612 1137 678
rect 1154 668 1158 671
rect 1146 658 1150 661
rect 1158 651 1161 658
rect 1150 648 1161 651
rect 1182 652 1185 738
rect 1278 722 1281 738
rect 1150 642 1153 648
rect 1182 632 1185 648
rect 898 568 902 571
rect 814 542 817 548
rect 774 482 777 488
rect 758 392 761 458
rect 758 352 761 388
rect 798 382 801 518
rect 838 492 841 548
rect 854 482 857 538
rect 822 472 825 478
rect 818 458 822 461
rect 862 452 865 458
rect 814 392 817 448
rect 782 362 785 368
rect 630 332 633 338
rect 670 332 673 338
rect 654 252 657 259
rect 670 192 673 268
rect 678 192 681 318
rect 686 262 689 268
rect 702 262 705 348
rect 722 338 726 341
rect 718 292 721 338
rect 578 168 582 171
rect 586 158 590 161
rect 522 148 526 151
rect 546 148 550 151
rect 518 132 521 138
rect 502 92 505 118
rect 534 82 537 138
rect 454 68 465 71
rect 366 62 369 68
rect 454 62 457 68
rect 418 58 422 61
rect 466 58 470 61
rect 254 52 257 58
rect 246 42 249 48
rect 270 -22 273 58
rect 446 52 449 58
rect 290 38 294 41
rect 476 3 477 7
rect 481 3 482 7
rect 486 3 488 7
rect 510 -19 513 68
rect 534 62 537 78
rect 542 72 545 148
rect 550 132 553 138
rect 558 102 561 148
rect 574 142 577 148
rect 598 132 601 148
rect 574 92 577 128
rect 582 82 585 108
rect 590 92 593 98
rect 554 78 558 81
rect 522 58 526 61
rect 554 58 558 61
rect 606 52 609 168
rect 678 162 681 168
rect 630 122 633 148
rect 646 142 649 148
rect 686 142 689 258
rect 702 142 705 258
rect 714 148 718 151
rect 642 138 646 141
rect 722 138 726 141
rect 642 128 646 131
rect 638 82 641 128
rect 670 72 673 138
rect 734 132 737 298
rect 750 282 753 318
rect 750 272 753 278
rect 782 272 785 358
rect 798 342 801 378
rect 846 342 849 368
rect 854 342 857 418
rect 870 392 873 438
rect 910 352 913 588
rect 938 548 942 551
rect 966 542 969 608
rect 974 552 977 598
rect 1078 582 1081 588
rect 1150 572 1153 578
rect 1010 558 1014 561
rect 1026 558 1030 561
rect 974 542 977 548
rect 1014 542 1017 548
rect 1038 542 1041 568
rect 1054 542 1057 558
rect 1062 542 1065 558
rect 1086 542 1089 558
rect 1126 552 1129 568
rect 1166 562 1169 628
rect 1190 602 1193 678
rect 1238 672 1241 678
rect 1238 652 1241 658
rect 1254 622 1257 668
rect 1270 652 1273 659
rect 1278 612 1281 718
rect 1294 672 1297 738
rect 1370 718 1374 721
rect 1382 702 1385 748
rect 1302 682 1305 688
rect 1374 672 1377 678
rect 1178 558 1182 561
rect 1134 542 1137 548
rect 1158 542 1161 548
rect 946 538 950 541
rect 1054 532 1057 538
rect 1062 532 1065 538
rect 1158 522 1161 528
rect 946 518 950 521
rect 988 503 989 507
rect 993 503 994 507
rect 998 503 1000 507
rect 1030 502 1033 518
rect 1046 492 1049 518
rect 1018 488 1022 491
rect 974 472 977 478
rect 1046 472 1049 488
rect 1062 472 1065 498
rect 1082 478 1086 481
rect 1070 471 1073 478
rect 1070 468 1078 471
rect 990 452 993 468
rect 1050 458 1054 461
rect 942 442 945 448
rect 922 418 926 421
rect 906 348 910 351
rect 854 322 857 338
rect 902 292 905 338
rect 942 332 945 378
rect 950 352 953 358
rect 970 348 974 351
rect 762 258 766 261
rect 822 252 825 278
rect 894 272 897 278
rect 834 258 838 261
rect 886 242 889 268
rect 690 128 694 131
rect 714 128 718 131
rect 718 92 721 108
rect 686 72 689 78
rect 734 72 737 118
rect 742 102 745 158
rect 798 142 801 238
rect 878 192 881 218
rect 866 188 870 191
rect 894 172 897 268
rect 926 262 929 318
rect 950 282 953 348
rect 998 342 1001 458
rect 1070 452 1073 458
rect 1014 362 1017 368
rect 958 272 961 318
rect 902 252 905 258
rect 942 252 945 268
rect 950 262 953 268
rect 966 262 969 338
rect 988 303 989 307
rect 993 303 994 307
rect 998 303 1000 307
rect 1014 292 1017 348
rect 1022 292 1025 398
rect 1034 358 1038 361
rect 1054 352 1057 358
rect 1070 352 1073 358
rect 1038 342 1041 348
rect 1078 342 1081 368
rect 1086 352 1089 448
rect 1094 432 1097 518
rect 1114 478 1118 481
rect 1134 472 1137 518
rect 1166 482 1169 558
rect 1174 542 1177 548
rect 1102 452 1105 468
rect 1110 452 1113 468
rect 1122 458 1126 461
rect 1134 442 1137 468
rect 1142 452 1145 468
rect 1158 452 1161 458
rect 1166 432 1169 468
rect 1174 452 1177 488
rect 1182 482 1185 558
rect 1190 552 1193 598
rect 1198 542 1201 608
rect 1234 558 1238 561
rect 1286 551 1289 558
rect 1254 542 1257 548
rect 1294 542 1297 668
rect 1358 662 1361 668
rect 1374 592 1377 618
rect 1382 542 1385 548
rect 1202 538 1206 541
rect 1254 532 1257 538
rect 1314 528 1318 531
rect 1222 462 1225 488
rect 1302 482 1305 498
rect 1186 458 1190 461
rect 1230 452 1233 478
rect 1254 462 1257 478
rect 1270 472 1273 478
rect 1358 472 1361 498
rect 1390 482 1393 668
rect 1398 592 1401 678
rect 1414 602 1417 658
rect 1422 592 1425 598
rect 1454 592 1457 808
rect 1446 582 1449 588
rect 1406 552 1409 568
rect 1282 468 1286 471
rect 1306 468 1310 471
rect 1186 438 1190 441
rect 1210 438 1214 441
rect 1102 342 1105 368
rect 1110 352 1113 418
rect 1126 362 1129 408
rect 1182 372 1185 418
rect 1210 358 1214 361
rect 1114 348 1118 351
rect 1182 342 1185 348
rect 1046 332 1049 338
rect 1066 328 1070 331
rect 1098 328 1102 331
rect 1146 318 1150 321
rect 1046 292 1049 308
rect 986 288 990 291
rect 990 252 993 258
rect 918 222 921 248
rect 982 242 985 248
rect 926 172 929 218
rect 942 192 945 238
rect 974 172 977 178
rect 962 168 966 171
rect 742 72 745 98
rect 798 92 801 138
rect 806 112 809 148
rect 846 91 849 148
rect 870 142 873 168
rect 890 158 894 161
rect 1010 158 1014 161
rect 1014 152 1017 158
rect 1022 152 1025 258
rect 1030 192 1033 258
rect 1054 252 1057 278
rect 1062 262 1065 268
rect 1070 242 1073 288
rect 1094 282 1097 318
rect 1158 282 1161 328
rect 1138 278 1142 281
rect 1086 272 1089 278
rect 1094 262 1097 278
rect 1102 262 1105 268
rect 1150 262 1153 278
rect 994 148 998 151
rect 902 132 905 148
rect 918 142 921 148
rect 862 122 865 128
rect 838 88 849 91
rect 838 82 841 88
rect 850 78 854 81
rect 806 72 809 78
rect 862 72 865 98
rect 870 92 873 108
rect 878 72 881 118
rect 886 82 889 118
rect 894 92 897 128
rect 910 112 913 138
rect 918 92 921 138
rect 974 102 977 148
rect 1030 122 1033 138
rect 1038 132 1041 168
rect 1062 122 1065 218
rect 1070 162 1073 168
rect 1078 152 1081 258
rect 1110 252 1113 258
rect 1130 238 1134 241
rect 1110 182 1113 218
rect 1086 142 1089 148
rect 1078 131 1081 138
rect 1094 131 1097 138
rect 1078 128 1097 131
rect 1102 132 1105 158
rect 1126 152 1129 158
rect 1134 142 1137 148
rect 988 103 989 107
rect 993 103 994 107
rect 998 103 1000 107
rect 1006 82 1009 98
rect 1062 91 1065 118
rect 1054 88 1065 91
rect 1070 92 1073 98
rect 818 68 822 71
rect 914 68 918 71
rect 982 70 985 78
rect 830 62 833 68
rect 654 42 657 59
rect 750 52 753 58
rect 854 52 857 58
rect 862 52 865 68
rect 934 62 937 68
rect 942 62 945 68
rect 1010 68 1014 71
rect 1054 62 1057 88
rect 1066 78 1070 81
rect 1102 72 1105 98
rect 1110 92 1113 128
rect 1118 121 1121 138
rect 1126 132 1129 138
rect 1118 118 1126 121
rect 1134 102 1137 138
rect 1142 82 1145 228
rect 1150 172 1153 258
rect 1158 162 1161 278
rect 1166 152 1169 338
rect 1198 332 1201 358
rect 1222 352 1225 428
rect 1230 412 1233 448
rect 1254 442 1257 448
rect 1262 432 1265 468
rect 1290 458 1294 461
rect 1342 452 1345 458
rect 1282 448 1286 451
rect 1310 362 1313 378
rect 1242 358 1246 361
rect 1338 358 1342 361
rect 1358 361 1361 468
rect 1390 452 1393 459
rect 1374 392 1377 438
rect 1398 392 1401 488
rect 1422 392 1425 538
rect 1430 502 1433 548
rect 1446 392 1449 558
rect 1462 541 1465 618
rect 1470 552 1473 708
rect 1462 538 1473 541
rect 1454 492 1457 498
rect 1454 381 1457 478
rect 1446 378 1457 381
rect 1350 358 1361 361
rect 1310 352 1313 358
rect 1226 338 1230 341
rect 1206 332 1209 338
rect 1222 272 1225 338
rect 1238 302 1241 348
rect 1314 338 1318 341
rect 1246 312 1249 328
rect 1254 322 1257 338
rect 1230 292 1233 298
rect 1238 282 1241 298
rect 1278 282 1281 288
rect 1286 262 1289 318
rect 1310 271 1313 318
rect 1318 281 1321 308
rect 1326 292 1329 338
rect 1334 312 1337 318
rect 1342 302 1345 358
rect 1350 342 1353 358
rect 1430 352 1433 358
rect 1318 278 1326 281
rect 1310 268 1318 271
rect 1226 258 1230 261
rect 1174 242 1177 258
rect 1182 252 1185 258
rect 1190 232 1193 258
rect 1202 238 1206 241
rect 1290 238 1294 241
rect 1118 72 1121 78
rect 1066 68 1070 71
rect 1158 62 1161 148
rect 1190 141 1193 218
rect 1186 138 1193 141
rect 1198 132 1201 158
rect 1206 152 1209 168
rect 1214 122 1217 138
rect 1222 132 1225 138
rect 1230 132 1233 178
rect 1238 162 1241 168
rect 1246 142 1249 148
rect 1302 142 1305 228
rect 1358 172 1361 348
rect 1366 262 1369 268
rect 1338 148 1342 151
rect 1310 142 1313 148
rect 1358 142 1361 148
rect 1374 142 1377 268
rect 1382 252 1385 348
rect 1406 292 1409 348
rect 1446 292 1449 378
rect 1454 362 1457 368
rect 1462 351 1465 518
rect 1454 348 1465 351
rect 1470 352 1473 538
rect 1454 292 1457 348
rect 1418 288 1422 291
rect 1430 191 1433 258
rect 1422 188 1433 191
rect 1394 148 1398 151
rect 1254 132 1257 138
rect 1302 132 1305 138
rect 1422 132 1425 188
rect 1442 138 1446 141
rect 1190 102 1193 118
rect 918 52 921 58
rect 1054 52 1057 58
rect 1078 52 1081 58
rect 1126 52 1129 58
rect 1174 52 1177 98
rect 1230 72 1233 118
rect 1246 72 1249 88
rect 1286 62 1289 118
rect 1326 92 1329 118
rect 1342 72 1345 88
rect 1390 72 1393 128
rect 1422 92 1425 128
rect 1358 63 1361 68
rect 1230 52 1233 58
rect 1262 52 1265 59
rect 1430 62 1433 108
rect 1446 92 1449 128
rect 1454 92 1457 278
rect 1478 262 1481 348
rect 1486 282 1489 378
rect 1470 62 1473 118
rect 1358 58 1361 59
rect 810 48 814 51
rect 942 42 945 48
rect 778 38 782 41
rect 510 -22 521 -19
rect 558 -22 561 8
<< m3contact >>
rect 158 1208 162 1212
rect 334 1208 338 1212
rect 230 1198 234 1202
rect 310 1198 314 1202
rect 190 1188 194 1192
rect 214 1178 218 1182
rect 238 1168 242 1172
rect 46 1148 50 1152
rect 366 1198 370 1202
rect 390 1198 394 1202
rect 382 1188 386 1192
rect 422 1188 426 1192
rect 430 1188 434 1192
rect 494 1208 498 1212
rect 472 1203 476 1207
rect 477 1203 481 1207
rect 482 1203 486 1207
rect 462 1198 466 1202
rect 454 1188 458 1192
rect 606 1208 610 1212
rect 646 1208 650 1212
rect 542 1198 546 1202
rect 566 1198 570 1202
rect 582 1198 586 1202
rect 526 1178 530 1182
rect 350 1158 354 1162
rect 366 1158 370 1162
rect 118 1148 122 1152
rect 206 1148 210 1152
rect 262 1148 266 1152
rect 286 1148 290 1152
rect 110 1128 114 1132
rect 94 1078 98 1082
rect 110 1078 114 1082
rect 54 1058 58 1062
rect 118 1058 122 1062
rect 134 1058 138 1062
rect 102 988 106 992
rect 54 948 58 952
rect 38 938 42 942
rect 118 938 122 942
rect 102 888 106 892
rect 190 1128 194 1132
rect 238 1138 242 1142
rect 214 1088 218 1092
rect 166 1078 170 1082
rect 174 1068 178 1072
rect 238 1068 242 1072
rect 182 968 186 972
rect 198 968 202 972
rect 166 958 170 962
rect 270 1138 274 1142
rect 294 1128 298 1132
rect 302 1128 306 1132
rect 318 1128 322 1132
rect 286 1118 290 1122
rect 270 1068 274 1072
rect 358 1068 362 1072
rect 350 1058 354 1062
rect 326 968 330 972
rect 222 948 226 952
rect 278 948 282 952
rect 142 888 146 892
rect 46 858 50 862
rect 118 858 122 862
rect 62 758 66 762
rect 230 878 234 882
rect 246 878 250 882
rect 270 878 274 882
rect 198 868 202 872
rect 310 888 314 892
rect 310 868 314 872
rect 182 858 186 862
rect 254 858 258 862
rect 294 858 298 862
rect 382 1108 386 1112
rect 398 1108 402 1112
rect 374 1098 378 1102
rect 694 1208 698 1212
rect 750 1208 754 1212
rect 686 1188 690 1192
rect 662 1178 666 1182
rect 734 1178 738 1182
rect 622 1168 626 1172
rect 630 1168 634 1172
rect 670 1168 674 1172
rect 686 1168 690 1172
rect 502 1158 506 1162
rect 630 1158 634 1162
rect 742 1158 746 1162
rect 438 1118 442 1122
rect 406 1088 410 1092
rect 422 1088 426 1092
rect 430 1058 434 1062
rect 398 968 402 972
rect 622 1148 626 1152
rect 478 1138 482 1142
rect 510 1138 514 1142
rect 478 1068 482 1072
rect 534 1068 538 1072
rect 566 1068 570 1072
rect 526 1048 530 1052
rect 534 1028 538 1032
rect 462 1018 466 1022
rect 454 978 458 982
rect 414 968 418 972
rect 430 968 434 972
rect 446 968 450 972
rect 398 948 402 952
rect 406 948 410 952
rect 382 928 386 932
rect 422 938 426 942
rect 446 948 450 952
rect 438 928 442 932
rect 398 888 402 892
rect 342 848 346 852
rect 366 848 370 852
rect 230 838 234 842
rect 206 818 210 822
rect 182 758 186 762
rect 198 758 202 762
rect 94 748 98 752
rect 174 748 178 752
rect 38 728 42 732
rect 6 688 10 692
rect 22 668 26 672
rect 30 658 34 662
rect 6 588 10 592
rect 30 558 34 562
rect 30 548 34 552
rect 54 548 58 552
rect 46 538 50 542
rect 54 518 58 522
rect 22 218 26 222
rect 150 738 154 742
rect 86 718 90 722
rect 102 718 106 722
rect 342 828 346 832
rect 222 748 226 752
rect 190 738 194 742
rect 190 718 194 722
rect 318 718 322 722
rect 262 708 266 712
rect 286 708 290 712
rect 318 708 322 712
rect 294 678 298 682
rect 238 668 242 672
rect 190 658 194 662
rect 238 658 242 662
rect 326 658 330 662
rect 374 808 378 812
rect 430 808 434 812
rect 422 778 426 782
rect 374 768 378 772
rect 358 658 362 662
rect 374 658 378 662
rect 374 648 378 652
rect 286 588 290 592
rect 230 578 234 582
rect 254 578 258 582
rect 302 578 306 582
rect 262 568 266 572
rect 70 558 74 562
rect 118 558 122 562
rect 206 558 210 562
rect 254 558 258 562
rect 86 548 90 552
rect 102 548 106 552
rect 174 548 178 552
rect 70 538 74 542
rect 86 528 90 532
rect 94 528 98 532
rect 118 528 122 532
rect 126 528 130 532
rect 102 488 106 492
rect 118 478 122 482
rect 54 398 58 402
rect 110 398 114 402
rect 110 388 114 392
rect 102 368 106 372
rect 110 368 114 372
rect 158 528 162 532
rect 166 518 170 522
rect 150 488 154 492
rect 142 468 146 472
rect 142 368 146 372
rect 126 358 130 362
rect 166 438 170 442
rect 158 358 162 362
rect 110 348 114 352
rect 134 348 138 352
rect 150 348 154 352
rect 86 338 90 342
rect 46 228 50 232
rect 38 218 42 222
rect 30 188 34 192
rect 14 158 18 162
rect 30 148 34 152
rect 70 318 74 322
rect 54 158 58 162
rect 62 158 66 162
rect 70 158 74 162
rect 102 328 106 332
rect 230 538 234 542
rect 190 498 194 502
rect 198 478 202 482
rect 190 468 194 472
rect 182 458 186 462
rect 278 528 282 532
rect 238 518 242 522
rect 270 518 274 522
rect 254 498 258 502
rect 230 468 234 472
rect 262 478 266 482
rect 214 458 218 462
rect 182 448 186 452
rect 198 448 202 452
rect 270 458 274 462
rect 222 448 226 452
rect 198 438 202 442
rect 254 438 258 442
rect 190 398 194 402
rect 134 268 138 272
rect 110 258 114 262
rect 126 238 130 242
rect 142 188 146 192
rect 142 178 146 182
rect 118 168 122 172
rect 134 168 138 172
rect 110 158 114 162
rect 62 128 66 132
rect 86 148 90 152
rect 54 68 58 72
rect 62 58 66 62
rect 134 148 138 152
rect 126 118 130 122
rect 166 328 170 332
rect 182 328 186 332
rect 182 318 186 322
rect 166 288 170 292
rect 230 428 234 432
rect 214 378 218 382
rect 294 488 298 492
rect 286 438 290 442
rect 294 368 298 372
rect 254 348 258 352
rect 246 338 250 342
rect 222 328 226 332
rect 246 328 250 332
rect 206 298 210 302
rect 158 268 162 272
rect 182 268 186 272
rect 166 248 170 252
rect 198 248 202 252
rect 174 228 178 232
rect 246 288 250 292
rect 222 278 226 282
rect 214 268 218 272
rect 254 278 258 282
rect 262 278 266 282
rect 414 728 418 732
rect 422 728 426 732
rect 398 668 402 672
rect 406 588 410 592
rect 472 1003 476 1007
rect 477 1003 481 1007
rect 482 1003 486 1007
rect 638 1138 642 1142
rect 622 1118 626 1122
rect 614 1108 618 1112
rect 582 1058 586 1062
rect 598 1058 602 1062
rect 574 998 578 1002
rect 622 1068 626 1072
rect 614 1048 618 1052
rect 630 1018 634 1022
rect 638 998 642 1002
rect 606 988 610 992
rect 566 968 570 972
rect 582 968 586 972
rect 478 958 482 962
rect 526 958 530 962
rect 534 958 538 962
rect 518 948 522 952
rect 526 938 530 942
rect 550 938 554 942
rect 494 928 498 932
rect 478 868 482 872
rect 566 878 570 882
rect 590 878 594 882
rect 526 868 530 872
rect 510 858 514 862
rect 550 848 554 852
rect 670 1118 674 1122
rect 798 1198 802 1202
rect 790 1178 794 1182
rect 758 1168 762 1172
rect 774 1168 778 1172
rect 766 1158 770 1162
rect 862 1178 866 1182
rect 862 1158 866 1162
rect 718 1138 722 1142
rect 766 1138 770 1142
rect 750 1108 754 1112
rect 686 1098 690 1102
rect 710 1098 714 1102
rect 814 1148 818 1152
rect 822 1148 826 1152
rect 798 1088 802 1092
rect 662 1068 666 1072
rect 902 1188 906 1192
rect 886 1138 890 1142
rect 1038 1208 1042 1212
rect 1022 1198 1026 1202
rect 982 1188 986 1192
rect 950 1178 954 1182
rect 966 1178 970 1182
rect 1046 1178 1050 1182
rect 942 1168 946 1172
rect 934 1148 938 1152
rect 982 1158 986 1162
rect 1038 1158 1042 1162
rect 966 1148 970 1152
rect 1030 1148 1034 1152
rect 846 1128 850 1132
rect 926 1128 930 1132
rect 942 1128 946 1132
rect 830 1118 834 1122
rect 926 1108 930 1112
rect 862 1098 866 1102
rect 894 1098 898 1102
rect 902 1098 906 1102
rect 838 1078 842 1082
rect 830 1068 834 1072
rect 782 1058 786 1062
rect 806 1058 810 1062
rect 654 1038 658 1042
rect 910 1078 914 1082
rect 854 1068 858 1072
rect 878 1068 882 1072
rect 742 1048 746 1052
rect 830 1048 834 1052
rect 790 1008 794 1012
rect 718 998 722 1002
rect 766 998 770 1002
rect 686 968 690 972
rect 670 938 674 942
rect 654 928 658 932
rect 638 868 642 872
rect 782 988 786 992
rect 718 958 722 962
rect 830 988 834 992
rect 830 968 834 972
rect 846 968 850 972
rect 846 958 850 962
rect 742 948 746 952
rect 790 948 794 952
rect 822 948 826 952
rect 702 938 706 942
rect 718 938 722 942
rect 734 938 738 942
rect 686 888 690 892
rect 726 928 730 932
rect 782 938 786 942
rect 750 908 754 912
rect 718 898 722 902
rect 798 938 802 942
rect 798 928 802 932
rect 862 938 866 942
rect 822 928 826 932
rect 814 918 818 922
rect 814 888 818 892
rect 734 878 738 882
rect 798 878 802 882
rect 710 868 714 872
rect 750 868 754 872
rect 614 858 618 862
rect 726 858 730 862
rect 606 828 610 832
rect 510 808 514 812
rect 472 803 476 807
rect 477 803 481 807
rect 482 803 486 807
rect 486 778 490 782
rect 502 758 506 762
rect 454 748 458 752
rect 438 738 442 742
rect 478 728 482 732
rect 622 818 626 822
rect 646 818 650 822
rect 622 798 626 802
rect 550 768 554 772
rect 558 768 562 772
rect 614 768 618 772
rect 574 758 578 762
rect 518 738 522 742
rect 502 708 506 712
rect 430 658 434 662
rect 422 638 426 642
rect 414 578 418 582
rect 390 568 394 572
rect 318 558 322 562
rect 358 558 362 562
rect 334 538 338 542
rect 382 548 386 552
rect 422 538 426 542
rect 350 518 354 522
rect 358 478 362 482
rect 318 448 322 452
rect 334 448 338 452
rect 334 438 338 442
rect 326 428 330 432
rect 310 398 314 402
rect 302 338 306 342
rect 294 328 298 332
rect 310 328 314 332
rect 278 308 282 312
rect 238 268 242 272
rect 286 298 290 302
rect 302 278 306 282
rect 230 258 234 262
rect 270 258 274 262
rect 214 248 218 252
rect 238 188 242 192
rect 158 178 162 182
rect 174 178 178 182
rect 166 148 170 152
rect 166 138 170 142
rect 150 108 154 112
rect 214 178 218 182
rect 230 168 234 172
rect 238 168 242 172
rect 214 148 218 152
rect 222 148 226 152
rect 198 118 202 122
rect 182 98 186 102
rect 198 88 202 92
rect 190 78 194 82
rect 206 78 210 82
rect 254 238 258 242
rect 278 238 282 242
rect 246 138 250 142
rect 238 118 242 122
rect 286 188 290 192
rect 318 318 322 322
rect 414 528 418 532
rect 398 518 402 522
rect 454 648 458 652
rect 472 603 476 607
rect 477 603 481 607
rect 482 603 486 607
rect 526 718 530 722
rect 510 698 514 702
rect 518 698 522 702
rect 742 798 746 802
rect 630 768 634 772
rect 646 758 650 762
rect 686 758 690 762
rect 702 758 706 762
rect 598 748 602 752
rect 574 738 578 742
rect 582 738 586 742
rect 614 738 618 742
rect 638 738 642 742
rect 646 738 650 742
rect 670 738 674 742
rect 542 728 546 732
rect 566 728 570 732
rect 606 718 610 722
rect 614 708 618 712
rect 614 698 618 702
rect 630 678 634 682
rect 566 668 570 672
rect 598 668 602 672
rect 558 658 562 662
rect 590 658 594 662
rect 606 658 610 662
rect 790 848 794 852
rect 814 848 818 852
rect 846 918 850 922
rect 782 838 786 842
rect 766 808 770 812
rect 758 768 762 772
rect 766 768 770 772
rect 718 728 722 732
rect 726 698 730 702
rect 662 678 666 682
rect 750 708 754 712
rect 758 698 762 702
rect 918 1058 922 1062
rect 902 1048 906 1052
rect 926 1038 930 1042
rect 942 1038 946 1042
rect 984 1103 988 1107
rect 989 1103 993 1107
rect 994 1103 998 1107
rect 1014 1128 1018 1132
rect 966 1048 970 1052
rect 958 1038 962 1042
rect 950 1018 954 1022
rect 926 1008 930 1012
rect 958 968 962 972
rect 1022 1098 1026 1102
rect 1038 1088 1042 1092
rect 1038 1078 1042 1082
rect 1078 1208 1082 1212
rect 1054 1168 1058 1172
rect 1062 1168 1066 1172
rect 1118 1208 1122 1212
rect 1110 1198 1114 1202
rect 1102 1188 1106 1192
rect 1150 1188 1154 1192
rect 1142 1178 1146 1182
rect 1198 1208 1202 1212
rect 1182 1198 1186 1202
rect 1238 1198 1242 1202
rect 1166 1178 1170 1182
rect 1206 1178 1210 1182
rect 1222 1178 1226 1182
rect 1222 1168 1226 1172
rect 1174 1158 1178 1162
rect 1086 1148 1090 1152
rect 1126 1148 1130 1152
rect 1134 1148 1138 1152
rect 1222 1148 1226 1152
rect 1246 1148 1250 1152
rect 1078 1138 1082 1142
rect 1102 1138 1106 1142
rect 1126 1138 1130 1142
rect 1158 1138 1162 1142
rect 1054 1098 1058 1102
rect 1070 1078 1074 1082
rect 1102 1118 1106 1122
rect 1142 1108 1146 1112
rect 1142 1098 1146 1102
rect 1134 1088 1138 1092
rect 1062 1068 1066 1072
rect 1078 1068 1082 1072
rect 1014 1058 1018 1062
rect 1030 1058 1034 1062
rect 1006 1048 1010 1052
rect 1070 1048 1074 1052
rect 1094 1058 1098 1062
rect 1118 1078 1122 1082
rect 1166 1068 1170 1072
rect 1278 1208 1282 1212
rect 1286 1198 1290 1202
rect 1270 1188 1274 1192
rect 1262 1138 1266 1142
rect 1190 1128 1194 1132
rect 1214 1088 1218 1092
rect 1206 1078 1210 1082
rect 1174 1058 1178 1062
rect 1190 1058 1194 1062
rect 1086 1038 1090 1042
rect 1030 1018 1034 1022
rect 910 948 914 952
rect 878 908 882 912
rect 886 888 890 892
rect 870 858 874 862
rect 862 828 866 832
rect 838 808 842 812
rect 822 798 826 802
rect 814 778 818 782
rect 806 768 810 772
rect 806 758 810 762
rect 870 798 874 802
rect 918 918 922 922
rect 958 918 962 922
rect 990 918 994 922
rect 942 908 946 912
rect 934 898 938 902
rect 918 878 922 882
rect 934 878 938 882
rect 942 858 946 862
rect 984 903 988 907
rect 989 903 993 907
rect 994 903 998 907
rect 974 878 978 882
rect 982 868 986 872
rect 966 858 970 862
rect 950 848 954 852
rect 966 848 970 852
rect 926 828 930 832
rect 918 818 922 822
rect 910 808 914 812
rect 902 778 906 782
rect 878 768 882 772
rect 894 768 898 772
rect 830 748 834 752
rect 822 738 826 742
rect 830 738 834 742
rect 782 728 786 732
rect 926 748 930 752
rect 862 738 866 742
rect 854 728 858 732
rect 902 718 906 722
rect 854 698 858 702
rect 846 688 850 692
rect 798 678 802 682
rect 646 668 650 672
rect 686 668 690 672
rect 734 668 738 672
rect 750 668 754 672
rect 830 668 834 672
rect 638 648 642 652
rect 782 658 786 662
rect 862 678 866 682
rect 886 678 890 682
rect 910 678 914 682
rect 878 668 882 672
rect 702 648 706 652
rect 766 648 770 652
rect 670 638 674 642
rect 614 598 618 602
rect 638 598 642 602
rect 654 598 658 602
rect 486 588 490 592
rect 566 588 570 592
rect 614 588 618 592
rect 526 568 530 572
rect 582 558 586 562
rect 646 588 650 592
rect 454 538 458 542
rect 462 538 466 542
rect 446 528 450 532
rect 438 498 442 502
rect 446 478 450 482
rect 630 548 634 552
rect 830 638 834 642
rect 750 618 754 622
rect 726 588 730 592
rect 686 568 690 572
rect 702 568 706 572
rect 678 548 682 552
rect 718 548 722 552
rect 566 538 570 542
rect 614 538 618 542
rect 462 488 466 492
rect 542 488 546 492
rect 502 478 506 482
rect 382 468 386 472
rect 438 468 442 472
rect 510 468 514 472
rect 374 458 378 462
rect 382 448 386 452
rect 350 398 354 402
rect 382 368 386 372
rect 414 448 418 452
rect 454 448 458 452
rect 510 448 514 452
rect 558 448 562 452
rect 534 438 538 442
rect 558 438 562 442
rect 446 428 450 432
rect 472 403 476 407
rect 477 403 481 407
rect 482 403 486 407
rect 454 378 458 382
rect 406 368 410 372
rect 422 368 426 372
rect 398 358 402 362
rect 374 348 378 352
rect 350 338 354 342
rect 374 338 378 342
rect 350 318 354 322
rect 318 268 322 272
rect 310 258 314 262
rect 326 248 330 252
rect 278 178 282 182
rect 294 178 298 182
rect 270 168 274 172
rect 270 148 274 152
rect 270 138 274 142
rect 262 128 266 132
rect 246 78 250 82
rect 198 68 202 72
rect 198 58 202 62
rect 214 58 218 62
rect 94 48 98 52
rect 294 158 298 162
rect 414 318 418 322
rect 374 278 378 282
rect 398 278 402 282
rect 502 358 506 362
rect 486 348 490 352
rect 446 338 450 342
rect 422 268 426 272
rect 382 258 386 262
rect 446 258 450 262
rect 390 248 394 252
rect 350 188 354 192
rect 326 178 330 182
rect 342 178 346 182
rect 318 138 322 142
rect 342 168 346 172
rect 390 168 394 172
rect 446 178 450 182
rect 422 158 426 162
rect 454 158 458 162
rect 374 148 378 152
rect 406 148 410 152
rect 446 148 450 152
rect 526 288 530 292
rect 598 528 602 532
rect 574 478 578 482
rect 590 468 594 472
rect 606 458 610 462
rect 718 458 722 462
rect 670 448 674 452
rect 662 438 666 442
rect 574 388 578 392
rect 590 378 594 382
rect 638 378 642 382
rect 662 378 666 382
rect 630 368 634 372
rect 574 358 578 362
rect 630 358 634 362
rect 614 338 618 342
rect 574 328 578 332
rect 566 278 570 282
rect 534 268 538 272
rect 472 203 476 207
rect 477 203 481 207
rect 482 203 486 207
rect 558 258 562 262
rect 542 248 546 252
rect 510 238 514 242
rect 566 238 570 242
rect 486 178 490 182
rect 510 178 514 182
rect 470 158 474 162
rect 438 138 442 142
rect 454 138 458 142
rect 462 138 466 142
rect 342 128 346 132
rect 382 128 386 132
rect 318 98 322 102
rect 326 98 330 102
rect 310 88 314 92
rect 390 98 394 102
rect 334 88 338 92
rect 374 78 378 82
rect 398 88 402 92
rect 326 68 330 72
rect 350 68 354 72
rect 366 68 370 72
rect 494 168 498 172
rect 502 148 506 152
rect 598 308 602 312
rect 614 268 618 272
rect 598 248 602 252
rect 614 248 618 252
rect 582 188 586 192
rect 646 348 650 352
rect 678 418 682 422
rect 718 408 722 412
rect 710 368 714 372
rect 694 358 698 362
rect 942 738 946 742
rect 926 728 930 732
rect 934 698 938 702
rect 982 818 986 822
rect 1126 978 1130 982
rect 1046 958 1050 962
rect 1062 958 1066 962
rect 1142 958 1146 962
rect 1166 988 1170 992
rect 1110 948 1114 952
rect 1158 948 1162 952
rect 1022 928 1026 932
rect 1054 938 1058 942
rect 1078 938 1082 942
rect 1086 938 1090 942
rect 1030 918 1034 922
rect 1046 918 1050 922
rect 1054 918 1058 922
rect 1086 918 1090 922
rect 1046 898 1050 902
rect 1182 978 1186 982
rect 1198 968 1202 972
rect 1230 1058 1234 1062
rect 1262 1078 1266 1082
rect 1246 1058 1250 1062
rect 1294 1148 1298 1152
rect 1318 1208 1322 1212
rect 1350 1208 1354 1212
rect 1342 1198 1346 1202
rect 1326 1188 1330 1192
rect 1318 1148 1322 1152
rect 1342 1148 1346 1152
rect 1318 1138 1322 1142
rect 1214 1048 1218 1052
rect 1230 1048 1234 1052
rect 1278 1048 1282 1052
rect 1214 1028 1218 1032
rect 1366 1208 1370 1212
rect 1366 1178 1370 1182
rect 1358 1138 1362 1142
rect 1398 1208 1402 1212
rect 1438 1208 1442 1212
rect 1430 1198 1434 1202
rect 1502 1228 1506 1232
rect 1478 1208 1482 1212
rect 1462 1188 1466 1192
rect 1390 1178 1394 1182
rect 1438 1168 1442 1172
rect 1382 1158 1386 1162
rect 1382 1148 1386 1152
rect 1398 1148 1402 1152
rect 1414 1148 1418 1152
rect 1430 1148 1434 1152
rect 1374 1128 1378 1132
rect 1414 1138 1418 1142
rect 1358 1068 1362 1072
rect 1326 1058 1330 1062
rect 1342 1048 1346 1052
rect 1246 988 1250 992
rect 1222 968 1226 972
rect 1278 958 1282 962
rect 1398 1078 1402 1082
rect 1382 1048 1386 1052
rect 1478 1158 1482 1162
rect 1430 1058 1434 1062
rect 1446 1058 1450 1062
rect 1486 1058 1490 1062
rect 1438 1008 1442 1012
rect 1358 958 1362 962
rect 1438 958 1442 962
rect 1462 958 1466 962
rect 1262 948 1266 952
rect 1318 948 1322 952
rect 1326 948 1330 952
rect 1390 948 1394 952
rect 1406 948 1410 952
rect 1430 948 1434 952
rect 1158 928 1162 932
rect 1166 908 1170 912
rect 1102 898 1106 902
rect 1062 878 1066 882
rect 1094 878 1098 882
rect 1086 868 1090 872
rect 1134 868 1138 872
rect 1142 868 1146 872
rect 1158 868 1162 872
rect 1022 858 1026 862
rect 1070 848 1074 852
rect 1102 848 1106 852
rect 1054 838 1058 842
rect 1086 838 1090 842
rect 1086 818 1090 822
rect 1046 808 1050 812
rect 1030 798 1034 802
rect 1238 918 1242 922
rect 1198 898 1202 902
rect 1190 888 1194 892
rect 1182 878 1186 882
rect 1198 878 1202 882
rect 1174 868 1178 872
rect 1182 858 1186 862
rect 1222 868 1226 872
rect 1222 858 1226 862
rect 1246 868 1250 872
rect 1294 868 1298 872
rect 1310 868 1314 872
rect 1270 858 1274 862
rect 1278 848 1282 852
rect 1286 838 1290 842
rect 1238 818 1242 822
rect 1206 808 1210 812
rect 1062 768 1066 772
rect 1046 758 1050 762
rect 966 738 970 742
rect 1014 738 1018 742
rect 958 728 962 732
rect 1006 728 1010 732
rect 950 718 954 722
rect 998 718 1002 722
rect 1014 708 1018 712
rect 984 703 988 707
rect 989 703 993 707
rect 994 703 998 707
rect 966 688 970 692
rect 918 658 922 662
rect 1222 758 1226 762
rect 1182 748 1186 752
rect 1254 748 1258 752
rect 1342 858 1346 862
rect 1398 858 1402 862
rect 1382 818 1386 822
rect 1406 818 1410 822
rect 1398 798 1402 802
rect 1342 788 1346 792
rect 1422 788 1426 792
rect 1462 918 1466 922
rect 1486 898 1490 902
rect 1478 838 1482 842
rect 1454 808 1458 812
rect 1486 808 1490 812
rect 1062 738 1066 742
rect 1094 738 1098 742
rect 1182 738 1186 742
rect 1222 738 1226 742
rect 1310 738 1314 742
rect 1046 718 1050 722
rect 1158 708 1162 712
rect 1174 708 1178 712
rect 1086 698 1090 702
rect 1086 688 1090 692
rect 1086 678 1090 682
rect 1078 668 1082 672
rect 1110 668 1114 672
rect 1006 658 1010 662
rect 942 648 946 652
rect 1150 668 1154 672
rect 1142 658 1146 662
rect 1278 718 1282 722
rect 1190 678 1194 682
rect 1238 678 1242 682
rect 1166 628 1170 632
rect 1182 628 1186 632
rect 966 608 970 612
rect 1134 608 1138 612
rect 910 588 914 592
rect 950 588 954 592
rect 902 568 906 572
rect 814 548 818 552
rect 774 488 778 492
rect 742 448 746 452
rect 758 388 762 392
rect 838 488 842 492
rect 822 478 826 482
rect 814 458 818 462
rect 814 448 818 452
rect 862 448 866 452
rect 870 438 874 442
rect 854 418 858 422
rect 798 378 802 382
rect 782 368 786 372
rect 758 348 762 352
rect 630 338 634 342
rect 670 338 674 342
rect 670 268 674 272
rect 654 248 658 252
rect 686 268 690 272
rect 718 338 722 342
rect 734 298 738 302
rect 702 258 706 262
rect 678 188 682 192
rect 622 178 626 182
rect 582 168 586 172
rect 678 168 682 172
rect 582 158 586 162
rect 518 148 522 152
rect 550 148 554 152
rect 574 148 578 152
rect 534 138 538 142
rect 518 128 522 132
rect 502 118 506 122
rect 534 78 538 82
rect 254 58 258 62
rect 422 58 426 62
rect 462 58 466 62
rect 246 38 250 42
rect 446 48 450 52
rect 286 38 290 42
rect 472 3 476 7
rect 477 3 481 7
rect 482 3 486 7
rect 550 128 554 132
rect 574 128 578 132
rect 598 128 602 132
rect 558 98 562 102
rect 582 108 586 112
rect 590 98 594 102
rect 558 78 562 82
rect 542 68 546 72
rect 518 58 522 62
rect 550 58 554 62
rect 646 148 650 152
rect 710 148 714 152
rect 646 138 650 142
rect 670 138 674 142
rect 686 138 690 142
rect 718 138 722 142
rect 646 128 650 132
rect 630 118 634 122
rect 638 78 642 82
rect 846 368 850 372
rect 942 548 946 552
rect 974 598 978 602
rect 1078 588 1082 592
rect 1150 578 1154 582
rect 1038 568 1042 572
rect 1126 568 1130 572
rect 1014 558 1018 562
rect 1022 558 1026 562
rect 1014 548 1018 552
rect 1054 558 1058 562
rect 1062 558 1066 562
rect 1238 648 1242 652
rect 1270 648 1274 652
rect 1254 618 1258 622
rect 1366 718 1370 722
rect 1382 698 1386 702
rect 1302 688 1306 692
rect 1374 678 1378 682
rect 1398 678 1402 682
rect 1294 668 1298 672
rect 1198 608 1202 612
rect 1278 608 1282 612
rect 1190 598 1194 602
rect 1182 558 1186 562
rect 1134 548 1138 552
rect 950 538 954 542
rect 974 538 978 542
rect 1054 538 1058 542
rect 1086 538 1090 542
rect 1158 538 1162 542
rect 1062 528 1066 532
rect 1158 528 1162 532
rect 950 518 954 522
rect 1134 518 1138 522
rect 984 503 988 507
rect 989 503 993 507
rect 994 503 998 507
rect 1030 498 1034 502
rect 1062 498 1066 502
rect 1022 488 1026 492
rect 1046 488 1050 492
rect 974 478 978 482
rect 1070 478 1074 482
rect 1086 478 1090 482
rect 998 458 1002 462
rect 1046 458 1050 462
rect 990 448 994 452
rect 942 438 946 442
rect 926 418 930 422
rect 942 378 946 382
rect 902 348 906 352
rect 854 318 858 322
rect 950 358 954 362
rect 966 348 970 352
rect 902 288 906 292
rect 894 278 898 282
rect 750 268 754 272
rect 782 268 786 272
rect 766 258 770 262
rect 830 258 834 262
rect 822 248 826 252
rect 886 238 890 242
rect 742 158 746 162
rect 686 128 690 132
rect 710 128 714 132
rect 734 118 738 122
rect 718 108 722 112
rect 686 78 690 82
rect 878 218 882 222
rect 870 188 874 192
rect 1070 448 1074 452
rect 1022 398 1026 402
rect 1014 358 1018 362
rect 966 338 970 342
rect 998 338 1002 342
rect 950 278 954 282
rect 950 268 954 272
rect 926 258 930 262
rect 984 303 988 307
rect 989 303 993 307
rect 994 303 998 307
rect 1078 368 1082 372
rect 1038 358 1042 362
rect 1054 358 1058 362
rect 1070 358 1074 362
rect 1118 478 1122 482
rect 1174 538 1178 542
rect 1174 488 1178 492
rect 1166 478 1170 482
rect 1110 468 1114 472
rect 1118 458 1122 462
rect 1102 448 1106 452
rect 1142 448 1146 452
rect 1158 448 1162 452
rect 1134 438 1138 442
rect 1230 558 1234 562
rect 1286 558 1290 562
rect 1254 548 1258 552
rect 1358 658 1362 662
rect 1374 618 1378 622
rect 1206 538 1210 542
rect 1382 538 1386 542
rect 1222 528 1226 532
rect 1254 528 1258 532
rect 1310 528 1314 532
rect 1302 498 1306 502
rect 1358 498 1362 502
rect 1222 488 1226 492
rect 1182 478 1186 482
rect 1230 478 1234 482
rect 1254 478 1258 482
rect 1270 478 1274 482
rect 1190 458 1194 462
rect 1422 598 1426 602
rect 1470 708 1474 712
rect 1446 588 1450 592
rect 1406 568 1410 572
rect 1446 558 1450 562
rect 1422 538 1426 542
rect 1398 488 1402 492
rect 1278 468 1282 472
rect 1302 468 1306 472
rect 1182 438 1186 442
rect 1206 438 1210 442
rect 1094 428 1098 432
rect 1166 428 1170 432
rect 1222 428 1226 432
rect 1110 418 1114 422
rect 1102 368 1106 372
rect 1126 408 1130 412
rect 1182 368 1186 372
rect 1126 358 1130 362
rect 1214 358 1218 362
rect 1118 348 1122 352
rect 1038 338 1042 342
rect 1166 338 1170 342
rect 1182 338 1186 342
rect 1046 328 1050 332
rect 1070 328 1074 332
rect 1102 328 1106 332
rect 1158 328 1162 332
rect 1094 318 1098 322
rect 1142 318 1146 322
rect 1046 308 1050 312
rect 982 288 986 292
rect 1014 288 1018 292
rect 1070 288 1074 292
rect 1054 278 1058 282
rect 1022 258 1026 262
rect 902 248 906 252
rect 942 248 946 252
rect 990 248 994 252
rect 942 238 946 242
rect 982 238 986 242
rect 918 218 922 222
rect 870 168 874 172
rect 894 168 898 172
rect 926 168 930 172
rect 958 168 962 172
rect 974 168 978 172
rect 846 148 850 152
rect 742 98 746 102
rect 806 108 810 112
rect 798 88 802 92
rect 894 158 898 162
rect 1014 158 1018 162
rect 1062 268 1066 272
rect 1086 278 1090 282
rect 1142 278 1146 282
rect 1158 278 1162 282
rect 1078 258 1082 262
rect 1102 258 1106 262
rect 1150 258 1154 262
rect 1030 188 1034 192
rect 1038 168 1042 172
rect 902 148 906 152
rect 990 148 994 152
rect 1014 148 1018 152
rect 918 138 922 142
rect 862 128 866 132
rect 894 128 898 132
rect 886 118 890 122
rect 870 108 874 112
rect 862 98 866 102
rect 806 78 810 82
rect 846 78 850 82
rect 910 108 914 112
rect 1070 168 1074 172
rect 1110 248 1114 252
rect 1134 238 1138 242
rect 1142 228 1146 232
rect 1110 178 1114 182
rect 1102 158 1106 162
rect 1126 158 1130 162
rect 1086 138 1090 142
rect 1094 138 1098 142
rect 1118 138 1122 142
rect 1134 138 1138 142
rect 1030 118 1034 122
rect 1062 118 1066 122
rect 984 103 988 107
rect 989 103 993 107
rect 994 103 998 107
rect 974 98 978 102
rect 1006 98 1010 102
rect 1070 98 1074 102
rect 1102 98 1106 102
rect 982 78 986 82
rect 822 68 826 72
rect 862 68 866 72
rect 918 68 922 72
rect 942 68 946 72
rect 606 48 610 52
rect 750 58 754 62
rect 830 58 834 62
rect 1006 68 1010 72
rect 1070 78 1074 82
rect 1126 128 1130 132
rect 1134 98 1138 102
rect 1150 168 1154 172
rect 1158 158 1162 162
rect 1254 438 1258 442
rect 1294 458 1298 462
rect 1278 448 1282 452
rect 1342 448 1346 452
rect 1262 428 1266 432
rect 1230 408 1234 412
rect 1310 378 1314 382
rect 1246 358 1250 362
rect 1342 358 1346 362
rect 1390 448 1394 452
rect 1374 438 1378 442
rect 1430 498 1434 502
rect 1462 518 1466 522
rect 1454 498 1458 502
rect 1454 478 1458 482
rect 1430 358 1434 362
rect 1238 348 1242 352
rect 1310 348 1314 352
rect 1230 338 1234 342
rect 1206 328 1210 332
rect 1318 338 1322 342
rect 1326 338 1330 342
rect 1254 318 1258 322
rect 1246 308 1250 312
rect 1230 298 1234 302
rect 1238 298 1242 302
rect 1278 288 1282 292
rect 1318 308 1322 312
rect 1334 308 1338 312
rect 1342 298 1346 302
rect 1326 288 1330 292
rect 1222 258 1226 262
rect 1286 258 1290 262
rect 1182 248 1186 252
rect 1174 238 1178 242
rect 1206 238 1210 242
rect 1294 238 1298 242
rect 1190 228 1194 232
rect 1302 228 1306 232
rect 1142 78 1146 82
rect 1070 68 1074 72
rect 1118 68 1122 72
rect 1182 138 1186 142
rect 1230 178 1234 182
rect 1206 168 1210 172
rect 1198 158 1202 162
rect 1238 168 1242 172
rect 1246 148 1250 152
rect 1366 268 1370 272
rect 1358 168 1362 172
rect 1310 148 1314 152
rect 1334 148 1338 152
rect 1358 148 1362 152
rect 1454 358 1458 362
rect 1486 378 1490 382
rect 1478 348 1482 352
rect 1406 288 1410 292
rect 1414 288 1418 292
rect 1454 278 1458 282
rect 1382 248 1386 252
rect 1398 148 1402 152
rect 1446 138 1450 142
rect 1222 128 1226 132
rect 1254 128 1258 132
rect 1302 128 1306 132
rect 1422 128 1426 132
rect 1446 128 1450 132
rect 1214 118 1218 122
rect 1230 118 1234 122
rect 1326 118 1330 122
rect 1174 98 1178 102
rect 1190 98 1194 102
rect 934 58 938 62
rect 1078 58 1082 62
rect 1158 58 1162 62
rect 1246 88 1250 92
rect 1230 68 1234 72
rect 1342 88 1346 92
rect 1430 108 1434 112
rect 1358 68 1362 72
rect 1286 58 1290 62
rect 1486 278 1490 282
rect 806 48 810 52
rect 854 48 858 52
rect 918 48 922 52
rect 942 48 946 52
rect 1054 48 1058 52
rect 1126 48 1130 52
rect 1230 48 1234 52
rect 1262 48 1266 52
rect 654 38 658 42
rect 782 38 786 42
rect 558 8 562 12
<< metal3 >>
rect 1498 1228 1502 1231
rect 162 1208 318 1211
rect 338 1208 462 1211
rect 498 1208 606 1211
rect 650 1208 694 1211
rect 754 1208 1038 1211
rect 1082 1208 1118 1211
rect 1162 1208 1198 1211
rect 1282 1208 1286 1211
rect 1322 1208 1326 1211
rect 1370 1208 1398 1211
rect 1442 1208 1478 1211
rect 486 1203 488 1207
rect 234 1198 294 1201
rect 314 1198 350 1201
rect 362 1198 366 1201
rect 394 1198 462 1201
rect 546 1198 550 1201
rect 562 1198 566 1201
rect 578 1198 582 1201
rect 802 1198 1022 1201
rect 1114 1198 1182 1201
rect 1242 1198 1286 1201
rect 1346 1198 1350 1201
rect 1382 1198 1430 1201
rect 182 1188 190 1191
rect 194 1188 382 1191
rect 418 1188 422 1191
rect 434 1188 441 1191
rect 450 1188 454 1191
rect 466 1188 686 1191
rect 906 1188 910 1191
rect 986 1188 1078 1191
rect 1106 1188 1150 1191
rect 1158 1188 1270 1191
rect 1318 1188 1326 1191
rect 1382 1191 1385 1198
rect 1330 1188 1385 1191
rect 1390 1188 1462 1191
rect 206 1178 214 1181
rect 218 1178 526 1181
rect 666 1178 689 1181
rect 686 1172 689 1178
rect 866 1178 950 1181
rect 970 1178 1046 1181
rect 1158 1181 1161 1188
rect 1390 1182 1393 1188
rect 1146 1178 1161 1181
rect 1170 1178 1206 1181
rect 1226 1178 1366 1181
rect 242 1168 622 1171
rect 634 1168 670 1171
rect 734 1171 737 1178
rect 734 1168 758 1171
rect 790 1171 793 1178
rect 778 1168 793 1171
rect 946 1168 1054 1171
rect 1066 1168 1222 1171
rect 1346 1168 1438 1171
rect 354 1158 366 1161
rect 506 1158 630 1161
rect 634 1158 742 1161
rect 770 1158 862 1161
rect 874 1158 982 1161
rect 1042 1158 1174 1161
rect 1386 1158 1478 1161
rect 50 1148 118 1151
rect 210 1148 262 1151
rect 266 1148 286 1151
rect 626 1148 814 1151
rect 826 1148 934 1151
rect 970 1148 1030 1151
rect 1090 1148 1126 1151
rect 1138 1148 1222 1151
rect 1226 1148 1246 1151
rect 1298 1148 1318 1151
rect 1322 1148 1342 1151
rect 1386 1148 1398 1151
rect 1402 1148 1414 1151
rect 1418 1148 1430 1151
rect 242 1138 270 1141
rect 450 1138 478 1141
rect 514 1138 521 1141
rect 642 1138 718 1141
rect 770 1138 849 1141
rect 890 1138 1070 1141
rect 1082 1138 1102 1141
rect 1106 1138 1126 1141
rect 1138 1138 1158 1141
rect 1266 1138 1318 1141
rect 1362 1138 1414 1141
rect 846 1132 849 1138
rect 114 1128 190 1131
rect 298 1128 302 1131
rect 306 1128 318 1131
rect 930 1128 942 1131
rect 1018 1128 1166 1131
rect 1170 1128 1190 1131
rect 1322 1128 1374 1131
rect 290 1118 438 1121
rect 626 1118 670 1121
rect 834 1118 929 1121
rect 938 1118 1102 1121
rect 926 1112 929 1118
rect 386 1108 398 1111
rect 618 1108 750 1111
rect 1018 1108 1142 1111
rect 998 1103 1000 1107
rect 378 1098 406 1101
rect 690 1098 710 1101
rect 866 1098 894 1101
rect 906 1098 934 1101
rect 1026 1098 1054 1101
rect 1082 1098 1142 1101
rect 98 1088 214 1091
rect 410 1088 422 1091
rect 802 1088 913 1091
rect 1042 1088 1134 1091
rect 1218 1088 1222 1091
rect 910 1082 913 1088
rect 98 1078 110 1081
rect 114 1078 166 1081
rect 842 1078 870 1081
rect 914 1078 1038 1081
rect 1050 1078 1070 1081
rect 1082 1078 1118 1081
rect 1210 1078 1262 1081
rect 1282 1078 1398 1081
rect 178 1068 238 1071
rect 482 1068 534 1071
rect 538 1068 566 1071
rect 570 1068 622 1071
rect 626 1068 662 1071
rect 834 1068 854 1071
rect 882 1068 1062 1071
rect 1066 1068 1078 1071
rect 1170 1068 1233 1071
rect 1242 1068 1249 1071
rect 58 1058 118 1061
rect 174 1061 177 1068
rect 138 1058 177 1061
rect 270 1061 273 1068
rect 270 1058 350 1061
rect 358 1061 361 1068
rect 1230 1062 1233 1068
rect 1246 1062 1249 1068
rect 358 1058 430 1061
rect 546 1058 582 1061
rect 602 1058 638 1061
rect 642 1058 782 1061
rect 786 1058 806 1061
rect 810 1058 918 1061
rect 922 1058 1014 1061
rect 1018 1058 1030 1061
rect 1070 1058 1094 1061
rect 1178 1058 1190 1061
rect 1358 1061 1361 1068
rect 1330 1058 1361 1061
rect 1434 1058 1446 1061
rect 1490 1058 1513 1061
rect 1070 1052 1073 1058
rect 530 1048 614 1051
rect 654 1048 742 1051
rect 834 1048 902 1051
rect 906 1048 966 1051
rect 1002 1048 1006 1051
rect 1218 1048 1230 1051
rect 1282 1048 1342 1051
rect 1346 1048 1382 1051
rect 654 1042 657 1048
rect 930 1038 934 1041
rect 946 1038 950 1041
rect 954 1038 958 1041
rect 962 1038 1086 1041
rect 538 1028 1214 1031
rect 466 1018 630 1021
rect 634 1018 942 1021
rect 954 1018 1030 1021
rect 498 1008 790 1011
rect 930 1008 1438 1011
rect 486 1003 488 1007
rect 578 998 638 1001
rect 642 998 718 1001
rect 770 998 1046 1001
rect 1166 992 1169 998
rect 94 988 102 991
rect 610 988 782 991
rect 786 988 830 991
rect 1170 988 1246 991
rect 458 978 1006 981
rect 1130 978 1182 981
rect 186 968 198 971
rect 330 968 398 971
rect 418 968 430 971
rect 434 968 446 971
rect 570 968 582 971
rect 586 968 686 971
rect 834 968 846 971
rect 1074 968 1198 971
rect 1218 968 1222 971
rect 170 958 478 961
rect 482 958 526 961
rect 530 958 534 961
rect 722 958 846 961
rect 958 961 961 968
rect 958 958 1014 961
rect 1050 958 1062 961
rect 1146 958 1278 961
rect 1362 958 1438 961
rect 1442 958 1462 961
rect 58 948 222 951
rect 282 948 398 951
rect 402 948 406 951
rect 410 948 446 951
rect 522 948 534 951
rect 538 948 737 951
rect 746 948 790 951
rect 826 948 865 951
rect 914 948 1110 951
rect 1162 948 1262 951
rect 1322 948 1326 951
rect 1330 948 1390 951
rect 1394 948 1406 951
rect 1410 948 1430 951
rect 734 942 737 948
rect 862 942 865 948
rect 1054 942 1057 948
rect 42 938 118 941
rect 530 938 550 941
rect 554 938 670 941
rect 674 938 702 941
rect 706 938 718 941
rect 786 938 798 941
rect 1090 938 1161 941
rect 422 931 425 938
rect 386 928 425 931
rect 442 928 494 931
rect 658 928 726 931
rect 826 928 1022 931
rect 1078 931 1081 938
rect 1026 928 1081 931
rect 1158 932 1161 938
rect 798 921 801 928
rect 562 918 801 921
rect 818 918 846 921
rect 922 918 958 921
rect 978 918 990 921
rect 1034 918 1046 921
rect 1058 918 1086 921
rect 1090 918 1238 921
rect 1466 918 1513 921
rect 522 908 750 911
rect 754 908 878 911
rect 882 908 942 911
rect 1010 908 1166 911
rect 1170 908 1246 911
rect 998 903 1000 907
rect 722 898 934 901
rect 1050 898 1102 901
rect 1110 898 1198 901
rect 1490 898 1513 901
rect 106 888 142 891
rect 314 888 398 891
rect 402 888 409 891
rect 698 888 814 891
rect 818 888 886 891
rect 1110 891 1113 898
rect 890 888 1113 891
rect 1178 888 1190 891
rect 234 878 246 881
rect 250 878 270 881
rect 686 881 689 888
rect 974 882 977 888
rect 594 878 689 881
rect 738 878 798 881
rect 802 878 918 881
rect 926 878 934 881
rect 938 878 966 881
rect 1066 878 1094 881
rect 1202 878 1513 881
rect 202 868 310 871
rect 566 871 569 878
rect 530 868 638 871
rect 714 868 750 871
rect 754 868 982 871
rect 1062 871 1065 878
rect 1058 868 1065 871
rect 1090 868 1134 871
rect 1146 868 1153 871
rect 1162 868 1174 871
rect 1182 871 1185 878
rect 1182 868 1222 871
rect 1250 868 1294 871
rect 50 858 118 861
rect 186 858 254 861
rect 478 861 481 868
rect 298 858 345 861
rect 478 858 510 861
rect 618 858 726 861
rect 946 858 966 861
rect 1026 858 1142 861
rect 1174 858 1182 861
rect 1210 858 1222 861
rect 1310 861 1313 868
rect 1274 858 1313 861
rect 1346 858 1398 861
rect 1490 858 1513 861
rect 342 852 345 858
rect 370 848 462 851
rect 466 848 550 851
rect 642 848 790 851
rect 870 851 873 858
rect 818 848 873 851
rect 946 848 950 851
rect 970 848 1070 851
rect 1074 848 1102 851
rect 1106 848 1278 851
rect 234 838 566 841
rect 786 838 1054 841
rect 1090 838 1166 841
rect 1290 838 1478 841
rect 346 828 606 831
rect 866 828 926 831
rect 930 828 937 831
rect 210 818 622 821
rect 650 818 918 821
rect 986 818 1086 821
rect 1242 818 1382 821
rect 1386 818 1406 821
rect 378 808 430 811
rect 514 808 766 811
rect 842 808 910 811
rect 1050 808 1206 811
rect 1458 808 1486 811
rect 486 803 488 807
rect 626 798 694 801
rect 746 798 822 801
rect 826 798 870 801
rect 874 798 1030 801
rect 1402 798 1513 801
rect 402 788 1342 791
rect 426 778 486 781
rect 490 778 814 781
rect 1422 781 1425 788
rect 1422 778 1513 781
rect 378 768 550 771
rect 562 768 566 771
rect 618 768 630 771
rect 634 768 758 771
rect 770 768 806 771
rect 810 768 878 771
rect 902 771 905 778
rect 898 768 905 771
rect 66 758 182 761
rect 186 758 198 761
rect 506 758 574 761
rect 578 758 646 761
rect 650 758 686 761
rect 706 758 806 761
rect 810 758 926 761
rect 930 758 1046 761
rect 1062 761 1065 768
rect 1062 758 1070 761
rect 1226 758 1513 761
rect 454 752 457 758
rect 98 748 174 751
rect 178 748 222 751
rect 590 748 598 751
rect 602 748 822 751
rect 834 748 926 751
rect 930 748 1182 751
rect 1258 748 1313 751
rect 1310 742 1313 748
rect 154 738 190 741
rect 442 738 518 741
rect 522 738 574 741
rect 586 738 614 741
rect 618 738 638 741
rect 642 738 646 741
rect 650 738 670 741
rect 826 738 830 741
rect 926 738 942 741
rect 946 738 966 741
rect 970 738 1014 741
rect 1066 738 1094 741
rect 1186 738 1222 741
rect 42 728 193 731
rect 418 728 422 731
rect 426 728 478 731
rect 546 728 566 731
rect 722 728 782 731
rect 826 728 854 731
rect 862 731 865 738
rect 926 732 929 738
rect 862 728 894 731
rect 954 728 958 731
rect 962 728 1006 731
rect 190 722 193 728
rect 90 718 102 721
rect 322 718 526 721
rect 530 718 606 721
rect 906 718 950 721
rect 1002 718 1046 721
rect 1282 718 1366 721
rect 266 708 286 711
rect 290 708 318 711
rect 506 708 518 711
rect 618 708 750 711
rect 1018 708 1158 711
rect 1162 708 1174 711
rect 1178 708 1470 711
rect 998 703 1000 707
rect 514 698 518 701
rect 522 698 614 701
rect 730 698 758 701
rect 762 698 854 701
rect 858 698 934 701
rect 938 698 977 701
rect 1090 698 1382 701
rect 850 688 966 691
rect 974 691 977 698
rect 974 688 1086 691
rect 6 681 9 688
rect -26 678 9 681
rect 298 678 494 681
rect 634 678 662 681
rect 802 678 862 681
rect 890 678 910 681
rect 966 681 969 688
rect 966 678 1086 681
rect 1194 678 1238 681
rect 1302 681 1305 688
rect 1242 678 1305 681
rect 1402 678 1513 681
rect 26 668 238 671
rect 570 668 598 671
rect 602 668 646 671
rect 650 668 657 671
rect 690 668 734 671
rect 754 668 830 671
rect 882 668 1078 671
rect 1114 668 1150 671
rect 1374 671 1377 678
rect 1298 668 1377 671
rect -26 658 30 661
rect 194 658 238 661
rect 242 658 249 661
rect 330 658 358 661
rect 362 658 374 661
rect 398 661 401 668
rect 1006 662 1009 668
rect 398 658 406 661
rect 410 658 430 661
rect 454 658 462 661
rect 530 658 558 661
rect 562 658 590 661
rect 610 658 782 661
rect 786 658 918 661
rect 1146 658 1153 661
rect 1238 658 1273 661
rect 1362 658 1513 661
rect 454 652 457 658
rect 1238 652 1241 658
rect 1270 652 1273 658
rect 378 648 446 651
rect 642 648 702 651
rect 770 648 942 651
rect 674 638 830 641
rect 422 631 425 638
rect 422 628 1158 631
rect 1170 628 1182 631
rect 754 618 1254 621
rect 1378 618 1513 621
rect 970 608 1134 611
rect 1138 608 1198 611
rect 1202 608 1278 611
rect 486 603 488 607
rect 618 598 638 601
rect 642 598 654 601
rect 978 598 1190 601
rect 1426 598 1513 601
rect 290 588 406 591
rect 490 588 566 591
rect 570 588 614 591
rect 618 588 638 591
rect 650 588 726 591
rect 914 588 950 591
rect 6 581 9 588
rect -26 578 9 581
rect 258 578 302 581
rect 306 578 414 581
rect 1078 581 1081 588
rect 1078 578 1150 581
rect 1446 581 1449 588
rect 1446 578 1513 581
rect 230 571 233 578
rect 230 568 262 571
rect 394 568 526 571
rect 530 568 537 571
rect 906 568 1038 571
rect 1042 568 1126 571
rect 1130 568 1406 571
rect -26 558 30 561
rect 74 558 118 561
rect 122 558 182 561
rect 210 558 254 561
rect 266 558 318 561
rect 354 558 358 561
rect 686 561 689 568
rect 586 558 689 561
rect 702 561 705 568
rect 702 558 974 561
rect 1018 558 1022 561
rect 1026 558 1054 561
rect 1066 558 1182 561
rect 1234 558 1286 561
rect 1450 558 1513 561
rect 34 548 54 551
rect 90 548 97 551
rect 106 548 174 551
rect 178 548 382 551
rect 634 548 678 551
rect 946 548 1014 551
rect 1018 548 1134 551
rect 1138 548 1254 551
rect 50 538 70 541
rect 234 538 334 541
rect 338 538 422 541
rect 458 538 462 541
rect 466 538 566 541
rect 598 538 614 541
rect 718 541 721 548
rect 814 541 817 548
rect 618 538 817 541
rect 954 538 974 541
rect 1058 538 1086 541
rect 1162 538 1174 541
rect 1210 538 1382 541
rect 1426 538 1513 541
rect 598 532 601 538
rect 54 528 86 531
rect 90 528 94 531
rect 122 528 126 531
rect 130 528 158 531
rect 162 528 278 531
rect 282 528 414 531
rect 418 528 446 531
rect 954 528 1062 531
rect 1162 528 1222 531
rect 1258 528 1310 531
rect 1314 528 1321 531
rect 54 522 57 528
rect 170 518 230 521
rect 234 518 238 521
rect 354 518 398 521
rect 942 518 950 521
rect 954 518 1134 521
rect 1466 518 1513 521
rect 270 512 273 518
rect 998 503 1000 507
rect 194 498 254 501
rect 442 498 462 501
rect 1034 498 1062 501
rect 1306 498 1358 501
rect 1362 498 1430 501
rect 1434 498 1454 501
rect 106 488 150 491
rect 154 488 294 491
rect 298 488 462 491
rect 466 488 542 491
rect 842 488 1022 491
rect 1050 488 1174 491
rect 1178 488 1222 491
rect 1510 491 1513 501
rect 1402 488 1513 491
rect 202 478 262 481
rect 266 478 273 481
rect 362 478 446 481
rect 506 478 574 481
rect 774 481 777 488
rect 774 478 822 481
rect 826 478 950 481
rect 978 478 1070 481
rect 1090 478 1118 481
rect 1186 478 1230 481
rect 1234 478 1254 481
rect 1458 478 1513 481
rect 118 471 121 478
rect 118 468 142 471
rect 146 468 190 471
rect 194 468 230 471
rect 386 468 438 471
rect 442 468 510 471
rect 514 468 518 471
rect 594 468 1006 471
rect 1010 468 1110 471
rect 1166 471 1169 478
rect 1270 471 1273 478
rect 1114 468 1273 471
rect 1282 468 1302 471
rect 270 462 273 468
rect 186 458 214 461
rect 222 458 246 461
rect 378 458 417 461
rect 458 458 606 461
rect 610 458 718 461
rect 818 458 998 461
rect 1002 458 1046 461
rect 1050 458 1118 461
rect 1122 458 1150 461
rect 1158 458 1190 461
rect 1194 458 1294 461
rect 1342 458 1393 461
rect 1482 458 1513 461
rect 222 452 225 458
rect 414 452 417 458
rect 1158 452 1161 458
rect 1342 452 1345 458
rect 1390 452 1393 458
rect 186 448 198 451
rect 254 448 318 451
rect 338 448 382 451
rect 458 448 510 451
rect 514 448 558 451
rect 562 448 670 451
rect 746 448 814 451
rect 866 448 945 451
rect 994 448 1070 451
rect 1106 448 1142 451
rect 1254 448 1278 451
rect 254 442 257 448
rect 942 442 945 448
rect 1254 442 1257 448
rect 170 438 198 441
rect 290 438 334 441
rect 538 438 558 441
rect 666 438 870 441
rect 1138 438 1182 441
rect 1186 438 1206 441
rect 1378 438 1478 441
rect 1490 438 1513 441
rect 234 428 326 431
rect 1098 428 1166 431
rect 1170 428 1222 431
rect 1226 428 1262 431
rect 446 421 449 428
rect 446 418 678 421
rect 718 418 854 421
rect 930 418 1110 421
rect 1490 418 1513 421
rect 718 412 721 418
rect 1130 408 1230 411
rect 486 403 488 407
rect 58 398 110 401
rect 114 398 190 401
rect 194 398 310 401
rect 314 398 350 401
rect 1026 398 1513 401
rect 578 388 758 391
rect 110 381 113 388
rect 110 378 214 381
rect 234 378 454 381
rect 594 378 638 381
rect 642 378 662 381
rect 802 378 942 381
rect 946 378 1310 381
rect 1490 378 1513 381
rect 106 368 110 371
rect 114 368 142 371
rect 298 368 382 371
rect 410 368 422 371
rect 634 368 710 371
rect 850 368 1017 371
rect 1082 368 1102 371
rect 1106 368 1182 371
rect 130 358 158 361
rect 402 358 502 361
rect 578 358 630 361
rect 782 361 785 368
rect 1014 362 1017 368
rect 698 358 785 361
rect 1042 358 1054 361
rect 1074 358 1126 361
rect 1218 358 1246 361
rect 1346 358 1430 361
rect 1458 358 1513 361
rect 114 348 134 351
rect 138 348 150 351
rect 258 348 374 351
rect 522 348 646 351
rect 762 348 902 351
rect 950 351 953 358
rect 950 348 966 351
rect 1122 348 1238 351
rect 1314 348 1478 351
rect 90 338 238 341
rect 242 338 246 341
rect 306 338 350 341
rect 378 338 446 341
rect 486 341 489 348
rect 466 338 489 341
rect 618 338 630 341
rect 674 338 718 341
rect 970 338 998 341
rect 1002 338 1038 341
rect 1042 338 1166 341
rect 1170 338 1182 341
rect 1234 338 1318 341
rect 1322 338 1326 341
rect 106 328 166 331
rect 186 328 222 331
rect 250 328 294 331
rect 314 328 574 331
rect 1050 328 1054 331
rect 1074 328 1102 331
rect 1106 328 1158 331
rect 1178 328 1206 331
rect 74 318 182 321
rect 186 318 318 321
rect 354 318 414 321
rect 858 318 1094 321
rect 1146 318 1254 321
rect 282 308 598 311
rect 1050 308 1238 311
rect 1250 308 1318 311
rect 1322 308 1334 311
rect 998 303 1000 307
rect 210 298 286 301
rect 290 298 734 301
rect 1242 298 1342 301
rect 170 288 246 291
rect 258 288 526 291
rect 906 288 982 291
rect 1018 288 1070 291
rect 1230 291 1233 298
rect 1074 288 1233 291
rect 1266 288 1278 291
rect 1330 288 1406 291
rect 1410 288 1414 291
rect 226 278 254 281
rect 266 278 302 281
rect 306 278 374 281
rect 402 278 566 281
rect 954 278 1054 281
rect 1146 278 1158 281
rect 1458 278 1486 281
rect 138 268 142 271
rect 162 268 182 271
rect 210 268 214 271
rect 242 268 318 271
rect 426 268 534 271
rect 618 268 670 271
rect 690 268 750 271
rect 894 271 897 278
rect 786 268 897 271
rect 1086 271 1089 278
rect 1066 268 1089 271
rect 114 258 230 261
rect 250 258 270 261
rect 274 258 310 261
rect 386 258 446 261
rect 562 258 702 261
rect 770 258 830 261
rect 834 258 841 261
rect 950 261 953 268
rect 930 258 1022 261
rect 1026 258 1078 261
rect 1082 258 1102 261
rect 1106 258 1150 261
rect 1186 258 1222 261
rect 1366 261 1369 268
rect 1290 258 1369 261
rect 126 248 166 251
rect 170 248 190 251
rect 194 248 198 251
rect 218 248 326 251
rect 330 248 390 251
rect 546 248 598 251
rect 618 248 654 251
rect 826 248 902 251
rect 906 248 942 251
rect 946 248 990 251
rect 1114 248 1182 251
rect 1186 248 1382 251
rect 126 242 129 248
rect 258 238 278 241
rect 514 238 566 241
rect 890 238 942 241
rect 986 238 1134 241
rect 1178 238 1206 241
rect 1210 238 1294 241
rect 50 228 174 231
rect 1146 228 1190 231
rect 1194 228 1302 231
rect 26 218 38 221
rect 882 218 918 221
rect 486 203 488 207
rect 34 188 142 191
rect 226 188 238 191
rect 266 188 286 191
rect 290 188 350 191
rect 354 188 582 191
rect 602 188 678 191
rect 874 188 1030 191
rect 146 178 158 181
rect 178 178 214 181
rect 282 178 294 181
rect 330 178 342 181
rect 450 178 486 181
rect 490 178 510 181
rect 514 178 622 181
rect 1114 178 1230 181
rect 230 172 233 178
rect 238 172 241 178
rect 122 168 134 171
rect 138 168 230 171
rect 274 168 342 171
rect 394 168 486 171
rect 570 168 582 171
rect 586 168 678 171
rect 874 168 894 171
rect 930 168 958 171
rect 978 168 1038 171
rect 1154 168 1206 171
rect 18 158 54 161
rect 66 158 70 161
rect 74 158 110 161
rect 114 158 294 161
rect 298 158 422 161
rect 426 158 449 161
rect 458 158 470 161
rect 494 161 497 168
rect 474 158 497 161
rect 586 158 593 161
rect 746 158 894 161
rect 898 158 902 161
rect 1006 158 1014 161
rect 1070 161 1073 168
rect 1070 158 1102 161
rect 1130 158 1150 161
rect 1162 158 1198 161
rect 1238 161 1241 168
rect 1202 158 1241 161
rect 1358 162 1361 168
rect 446 152 449 158
rect 34 148 86 151
rect 138 148 166 151
rect 206 148 214 151
rect 226 148 270 151
rect 378 148 406 151
rect 506 148 518 151
rect 554 148 574 151
rect 650 148 710 151
rect 850 148 902 151
rect 906 148 990 151
rect 1018 148 1246 151
rect 1338 148 1342 151
rect 1386 148 1398 151
rect 170 138 246 141
rect 258 138 265 141
rect 274 138 318 141
rect 322 138 438 141
rect 442 138 454 141
rect 466 138 521 141
rect 538 138 646 141
rect 674 138 686 141
rect 722 138 729 141
rect 922 138 1086 141
rect 1098 138 1118 141
rect 1138 138 1182 141
rect 1222 138 1257 141
rect 1310 141 1313 148
rect 1306 138 1313 141
rect 1358 141 1361 148
rect 1358 138 1446 141
rect 262 132 265 138
rect 518 132 521 138
rect 550 132 553 138
rect 1222 132 1225 138
rect 1254 132 1257 138
rect 66 128 241 131
rect 346 128 382 131
rect 578 128 598 131
rect 650 128 686 131
rect 690 128 710 131
rect 898 128 1126 131
rect 1306 128 1422 131
rect 1450 128 1486 131
rect 238 122 241 128
rect 130 118 198 121
rect 506 118 630 121
rect 862 121 865 128
rect 738 118 886 121
rect 898 118 1009 121
rect 1034 118 1038 121
rect 1066 118 1214 121
rect 1234 118 1326 121
rect 1330 118 1358 121
rect 154 108 254 111
rect 586 108 598 111
rect 722 108 806 111
rect 874 108 910 111
rect 1006 111 1009 118
rect 1006 108 1430 111
rect 998 103 1000 107
rect 186 98 318 101
rect 330 98 390 101
rect 594 98 742 101
rect 866 98 974 101
rect 1010 98 1070 101
rect 1106 98 1134 101
rect 1178 98 1190 101
rect 558 92 561 98
rect 190 88 198 91
rect 202 88 310 91
rect 338 88 398 91
rect 802 88 1246 91
rect 1250 88 1342 91
rect 210 78 246 81
rect 258 78 374 81
rect 378 78 534 81
rect 562 78 638 81
rect 810 78 846 81
rect 986 78 1006 81
rect 1074 78 1142 81
rect 190 71 193 78
rect 58 68 193 71
rect 202 68 222 71
rect 330 68 350 71
rect 370 68 542 71
rect 686 71 689 78
rect 686 68 790 71
rect 826 68 862 71
rect 922 68 942 71
rect 946 68 1006 71
rect 1074 68 1118 71
rect 1122 68 1230 71
rect 66 58 198 61
rect 426 58 462 61
rect 522 58 550 61
rect 554 58 726 61
rect 834 58 934 61
rect 938 58 1078 61
rect 1082 58 1158 61
rect 1230 58 1265 61
rect 1358 61 1361 68
rect 1290 58 1361 61
rect 214 51 217 58
rect 254 51 257 58
rect 98 48 257 51
rect 450 48 606 51
rect 750 51 753 58
rect 1230 52 1233 58
rect 1262 52 1265 58
rect 750 48 806 51
rect 858 48 918 51
rect 1058 48 1126 51
rect 250 38 286 41
rect 658 38 782 41
rect 942 41 945 48
rect 794 38 945 41
rect 558 12 561 18
rect 486 3 488 7
<< m4contact >>
rect 1494 1228 1498 1232
rect 318 1208 322 1212
rect 462 1208 466 1212
rect 1158 1208 1162 1212
rect 1286 1208 1290 1212
rect 1326 1208 1330 1212
rect 1350 1208 1354 1212
rect 473 1203 476 1207
rect 476 1203 477 1207
rect 479 1203 481 1207
rect 481 1203 482 1207
rect 482 1203 483 1207
rect 294 1198 298 1202
rect 350 1198 354 1202
rect 358 1198 362 1202
rect 550 1198 554 1202
rect 558 1198 562 1202
rect 574 1198 578 1202
rect 1350 1198 1354 1202
rect 414 1188 418 1192
rect 430 1188 434 1192
rect 446 1188 450 1192
rect 462 1188 466 1192
rect 910 1188 914 1192
rect 1078 1188 1082 1192
rect 1342 1168 1346 1172
rect 870 1158 874 1162
rect 446 1138 450 1142
rect 510 1138 514 1142
rect 1070 1138 1074 1142
rect 1134 1138 1138 1142
rect 1166 1128 1170 1132
rect 1318 1128 1322 1132
rect 934 1118 938 1122
rect 926 1108 930 1112
rect 1014 1108 1018 1112
rect 985 1103 988 1107
rect 988 1103 989 1107
rect 991 1103 993 1107
rect 993 1103 994 1107
rect 994 1103 995 1107
rect 406 1098 410 1102
rect 934 1098 938 1102
rect 1078 1098 1082 1102
rect 94 1088 98 1092
rect 1222 1088 1226 1092
rect 870 1078 874 1082
rect 1046 1078 1050 1082
rect 1078 1078 1082 1082
rect 1278 1078 1282 1082
rect 1238 1068 1242 1072
rect 542 1058 546 1062
rect 638 1058 642 1062
rect 998 1048 1002 1052
rect 934 1038 938 1042
rect 950 1038 954 1042
rect 942 1018 946 1022
rect 494 1008 498 1012
rect 473 1003 476 1007
rect 476 1003 477 1007
rect 479 1003 481 1007
rect 481 1003 482 1007
rect 482 1003 483 1007
rect 1046 998 1050 1002
rect 1166 998 1170 1002
rect 102 988 106 992
rect 454 978 458 982
rect 1006 978 1010 982
rect 1070 968 1074 972
rect 1214 968 1218 972
rect 1014 958 1018 962
rect 534 948 538 952
rect 558 918 562 922
rect 974 918 978 922
rect 518 908 522 912
rect 1006 908 1010 912
rect 1246 908 1250 912
rect 985 903 988 907
rect 988 903 989 907
rect 991 903 993 907
rect 993 903 994 907
rect 994 903 995 907
rect 398 888 402 892
rect 694 888 698 892
rect 1174 888 1178 892
rect 966 878 970 882
rect 1054 868 1058 872
rect 1142 868 1146 872
rect 1142 858 1146 862
rect 1182 858 1186 862
rect 1206 858 1210 862
rect 1486 858 1490 862
rect 462 848 466 852
rect 638 848 642 852
rect 942 848 946 852
rect 566 838 570 842
rect 1166 838 1170 842
rect 473 803 476 807
rect 476 803 477 807
rect 479 803 481 807
rect 481 803 482 807
rect 482 803 483 807
rect 694 798 698 802
rect 398 788 402 792
rect 566 768 570 772
rect 454 758 458 762
rect 926 758 930 762
rect 1070 758 1074 762
rect 822 748 826 752
rect 822 728 826 732
rect 894 728 898 732
rect 950 728 954 732
rect 518 708 522 712
rect 985 703 988 707
rect 988 703 989 707
rect 991 703 993 707
rect 993 703 994 707
rect 994 703 995 707
rect 494 678 498 682
rect 406 658 410 662
rect 462 658 466 662
rect 526 658 530 662
rect 1142 658 1146 662
rect 446 648 450 652
rect 1158 628 1162 632
rect 473 603 476 607
rect 476 603 477 607
rect 479 603 481 607
rect 481 603 482 607
rect 482 603 483 607
rect 638 588 642 592
rect 182 558 186 562
rect 262 558 266 562
rect 350 558 354 562
rect 974 558 978 562
rect 86 548 90 552
rect 950 528 954 532
rect 230 518 234 522
rect 270 508 274 512
rect 985 503 988 507
rect 988 503 989 507
rect 991 503 993 507
rect 993 503 994 507
rect 994 503 995 507
rect 462 498 466 502
rect 950 478 954 482
rect 270 468 274 472
rect 518 468 522 472
rect 1006 468 1010 472
rect 246 458 250 462
rect 454 458 458 462
rect 1150 458 1154 462
rect 1478 458 1482 462
rect 1478 438 1482 442
rect 1486 438 1490 442
rect 1262 428 1266 432
rect 1486 418 1490 422
rect 473 403 476 407
rect 476 403 477 407
rect 479 403 481 407
rect 481 403 482 407
rect 482 403 483 407
rect 230 378 234 382
rect 1182 368 1186 372
rect 518 348 522 352
rect 238 338 242 342
rect 462 338 466 342
rect 574 328 578 332
rect 1054 328 1058 332
rect 1174 328 1178 332
rect 1238 308 1242 312
rect 985 303 988 307
rect 988 303 989 307
rect 991 303 993 307
rect 993 303 994 307
rect 994 303 995 307
rect 254 288 258 292
rect 1262 288 1266 292
rect 142 268 146 272
rect 206 268 210 272
rect 246 258 250 262
rect 1182 258 1186 262
rect 190 248 194 252
rect 473 203 476 207
rect 476 203 477 207
rect 479 203 481 207
rect 481 203 482 207
rect 482 203 483 207
rect 222 188 226 192
rect 262 188 266 192
rect 598 188 602 192
rect 230 178 234 182
rect 238 178 242 182
rect 486 168 490 172
rect 566 168 570 172
rect 582 158 586 162
rect 902 158 906 162
rect 1014 158 1018 162
rect 1150 158 1154 162
rect 1358 158 1362 162
rect 214 148 218 152
rect 1342 148 1346 152
rect 1382 148 1386 152
rect 254 138 258 142
rect 718 138 722 142
rect 1094 138 1098 142
rect 1302 138 1306 142
rect 1486 128 1490 132
rect 894 118 898 122
rect 1038 118 1042 122
rect 1358 118 1362 122
rect 254 108 258 112
rect 598 108 602 112
rect 985 103 988 107
rect 988 103 989 107
rect 991 103 993 107
rect 993 103 994 107
rect 994 103 995 107
rect 558 88 562 92
rect 190 78 194 82
rect 254 78 258 82
rect 1006 78 1010 82
rect 222 68 226 72
rect 790 68 794 72
rect 726 58 730 62
rect 790 38 794 42
rect 558 18 562 22
rect 473 3 476 7
rect 476 3 477 7
rect 479 3 481 7
rect 481 3 482 7
rect 482 3 483 7
<< metal4 >>
rect 1498 1228 1505 1231
rect 1502 1222 1505 1228
rect 322 1208 326 1211
rect 1278 1208 1286 1211
rect 1318 1208 1326 1211
rect 1354 1208 1358 1211
rect 298 1198 302 1201
rect 362 1198 369 1201
rect 350 1192 353 1198
rect 418 1188 425 1191
rect 434 1188 438 1191
rect 454 1191 457 1208
rect 450 1188 457 1191
rect 462 1192 465 1208
rect 486 1203 488 1207
rect 542 1198 550 1201
rect 562 1198 569 1201
rect 578 1198 585 1201
rect 514 1138 521 1141
rect 94 991 97 1088
rect 94 988 102 991
rect 406 891 409 1098
rect 402 888 409 891
rect 398 661 401 788
rect 398 658 406 661
rect 446 652 449 1138
rect 486 1003 488 1007
rect 454 762 457 978
rect 462 662 465 848
rect 486 803 488 807
rect 494 682 497 1008
rect 518 912 521 1138
rect 542 1062 545 1198
rect 526 948 534 951
rect 518 712 521 908
rect 526 662 529 948
rect 558 771 561 918
rect 566 842 569 1198
rect 582 1192 585 1198
rect 902 1188 910 1191
rect 870 1082 873 1158
rect 638 852 641 1058
rect 558 768 566 771
rect 454 658 462 661
rect 186 558 190 561
rect 354 558 361 561
rect 262 552 265 558
rect 90 548 102 551
rect 230 382 233 518
rect 270 472 273 508
rect 454 462 457 658
rect 486 603 488 607
rect 638 592 641 848
rect 694 802 697 888
rect 926 762 929 1108
rect 934 1102 937 1118
rect 998 1103 1000 1107
rect 1002 1048 1009 1051
rect 934 1042 937 1048
rect 942 1038 950 1041
rect 942 1022 945 1038
rect 942 852 945 1018
rect 966 872 969 878
rect 822 732 825 748
rect 898 728 902 731
rect 954 728 961 731
rect 974 562 977 918
rect 1006 912 1009 978
rect 1014 962 1017 1108
rect 1070 1091 1073 1138
rect 1078 1102 1081 1188
rect 1134 1142 1137 1188
rect 1070 1088 1081 1091
rect 1078 1082 1081 1088
rect 1046 1002 1049 1078
rect 998 903 1000 907
rect 1058 868 1065 871
rect 1070 762 1073 968
rect 1146 868 1150 871
rect 1146 858 1150 861
rect 998 703 1000 707
rect 1146 658 1153 661
rect 134 268 142 271
rect 190 82 193 248
rect 206 151 209 268
rect 206 148 214 151
rect 222 72 225 188
rect 230 182 233 378
rect 238 182 241 338
rect 246 262 249 458
rect 462 342 465 498
rect 950 482 953 528
rect 998 503 1000 507
rect 486 403 488 407
rect 518 352 521 468
rect 254 272 257 288
rect 486 203 488 207
rect 262 141 265 188
rect 574 171 577 328
rect 998 303 1000 307
rect 570 168 577 171
rect 486 162 489 168
rect 586 158 593 161
rect 258 138 265 141
rect 598 112 601 188
rect 894 158 902 161
rect 1006 161 1009 468
rect 1150 462 1153 658
rect 1158 632 1161 1208
rect 1166 1002 1169 1128
rect 1166 842 1169 998
rect 1222 971 1225 1088
rect 1278 1082 1281 1208
rect 1318 1132 1321 1208
rect 1342 1198 1350 1201
rect 1342 1172 1345 1198
rect 1242 1068 1249 1071
rect 1218 968 1225 971
rect 1246 912 1249 1068
rect 1174 861 1177 888
rect 1174 858 1182 861
rect 1214 861 1217 868
rect 1210 858 1217 861
rect 1482 858 1486 861
rect 1478 442 1481 458
rect 1046 328 1054 331
rect 1170 328 1174 331
rect 1182 262 1185 368
rect 1238 312 1241 438
rect 1486 432 1489 438
rect 1262 292 1265 428
rect 1006 158 1014 161
rect 722 138 729 141
rect 254 82 257 108
rect 558 22 561 88
rect 726 62 729 138
rect 894 122 897 158
rect 998 103 1000 107
rect 1006 82 1009 158
rect 1150 142 1153 158
rect 1346 148 1350 151
rect 1306 138 1313 141
rect 1094 122 1097 138
rect 1358 122 1361 158
rect 1386 148 1393 151
rect 1486 132 1489 418
rect 1030 118 1038 121
rect 790 42 793 68
rect 486 3 488 7
<< m5contact >>
rect 1502 1218 1506 1222
rect 326 1208 330 1212
rect 454 1208 458 1212
rect 1358 1208 1362 1212
rect 302 1198 306 1202
rect 358 1198 362 1202
rect 350 1188 354 1192
rect 414 1188 418 1192
rect 438 1188 442 1192
rect 472 1203 473 1207
rect 473 1203 476 1207
rect 477 1203 479 1207
rect 479 1203 481 1207
rect 482 1203 483 1207
rect 483 1203 486 1207
rect 472 1003 473 1007
rect 473 1003 476 1007
rect 477 1003 479 1007
rect 479 1003 481 1007
rect 482 1003 483 1007
rect 483 1003 486 1007
rect 472 803 473 807
rect 473 803 476 807
rect 477 803 479 807
rect 479 803 481 807
rect 482 803 483 807
rect 483 803 486 807
rect 582 1188 586 1192
rect 910 1188 914 1192
rect 1134 1188 1138 1192
rect 190 558 194 562
rect 350 558 354 562
rect 102 548 106 552
rect 262 548 266 552
rect 472 603 473 607
rect 473 603 476 607
rect 477 603 479 607
rect 479 603 481 607
rect 482 603 483 607
rect 483 603 486 607
rect 984 1103 985 1107
rect 985 1103 988 1107
rect 989 1103 991 1107
rect 991 1103 993 1107
rect 994 1103 995 1107
rect 995 1103 998 1107
rect 934 1048 938 1052
rect 998 1048 1002 1052
rect 966 868 970 872
rect 902 728 906 732
rect 950 728 954 732
rect 984 903 985 907
rect 985 903 988 907
rect 989 903 991 907
rect 991 903 993 907
rect 994 903 995 907
rect 995 903 998 907
rect 1054 868 1058 872
rect 1150 868 1154 872
rect 1150 858 1154 862
rect 984 703 985 707
rect 985 703 988 707
rect 989 703 991 707
rect 991 703 993 707
rect 994 703 995 707
rect 995 703 998 707
rect 142 268 146 272
rect 984 503 985 507
rect 985 503 988 507
rect 989 503 991 507
rect 991 503 993 507
rect 994 503 995 507
rect 995 503 998 507
rect 472 403 473 407
rect 473 403 476 407
rect 477 403 479 407
rect 479 403 481 407
rect 482 403 483 407
rect 483 403 486 407
rect 254 268 258 272
rect 472 203 473 207
rect 473 203 476 207
rect 477 203 479 207
rect 479 203 481 207
rect 482 203 483 207
rect 483 203 486 207
rect 984 303 985 307
rect 985 303 988 307
rect 989 303 991 307
rect 991 303 993 307
rect 994 303 995 307
rect 995 303 998 307
rect 486 158 490 162
rect 582 158 586 162
rect 1214 868 1218 872
rect 1478 858 1482 862
rect 1238 438 1242 442
rect 1054 328 1058 332
rect 1166 328 1170 332
rect 1486 428 1490 432
rect 984 103 985 107
rect 985 103 988 107
rect 989 103 991 107
rect 991 103 993 107
rect 994 103 995 107
rect 995 103 998 107
rect 1350 148 1354 152
rect 1150 138 1154 142
rect 1302 138 1306 142
rect 1382 148 1386 152
rect 1038 118 1042 122
rect 1094 118 1098 122
rect 472 3 473 7
rect 473 3 476 7
rect 477 3 479 7
rect 479 3 481 7
rect 482 3 483 7
rect 483 3 486 7
<< metal5 >>
rect 330 1208 454 1211
rect 1502 1211 1505 1218
rect 1362 1208 1505 1211
rect 486 1203 488 1207
rect 472 1202 473 1203
rect 478 1202 480 1203
rect 485 1202 488 1203
rect 306 1198 358 1201
rect 354 1188 414 1191
rect 442 1188 582 1191
rect 914 1188 1134 1191
rect 998 1103 1000 1107
rect 984 1102 985 1103
rect 990 1102 992 1103
rect 997 1102 1000 1103
rect 938 1048 998 1051
rect 486 1003 488 1007
rect 472 1002 473 1003
rect 478 1002 480 1003
rect 485 1002 488 1003
rect 998 903 1000 907
rect 984 902 985 903
rect 990 902 992 903
rect 997 902 1000 903
rect 970 868 1054 871
rect 1154 868 1214 871
rect 1154 858 1478 861
rect 486 803 488 807
rect 472 802 473 803
rect 478 802 480 803
rect 485 802 488 803
rect 906 728 950 731
rect 998 703 1000 707
rect 984 702 985 703
rect 990 702 992 703
rect 997 702 1000 703
rect 486 603 488 607
rect 472 602 473 603
rect 478 602 480 603
rect 485 602 488 603
rect 194 558 350 561
rect 106 548 262 551
rect 998 503 1000 507
rect 984 502 985 503
rect 990 502 992 503
rect 997 502 1000 503
rect 1242 438 1489 441
rect 1486 432 1489 438
rect 486 403 488 407
rect 472 402 473 403
rect 478 402 480 403
rect 485 402 488 403
rect 1058 328 1166 331
rect 998 303 1000 307
rect 984 302 985 303
rect 990 302 992 303
rect 997 302 1000 303
rect 146 268 254 271
rect 486 203 488 207
rect 472 202 473 203
rect 478 202 480 203
rect 485 202 488 203
rect 490 158 582 161
rect 1354 148 1382 151
rect 1154 138 1302 141
rect 1042 118 1094 121
rect 998 103 1000 107
rect 984 102 985 103
rect 990 102 992 103
rect 997 102 1000 103
rect 486 3 488 7
rect 472 2 473 3
rect 478 2 480 3
rect 485 2 488 3
<< m6contact >>
rect 473 1203 476 1207
rect 476 1203 477 1207
rect 477 1203 478 1207
rect 480 1203 481 1207
rect 481 1203 482 1207
rect 482 1203 485 1207
rect 473 1202 478 1203
rect 480 1202 485 1203
rect 985 1103 988 1107
rect 988 1103 989 1107
rect 989 1103 990 1107
rect 992 1103 993 1107
rect 993 1103 994 1107
rect 994 1103 997 1107
rect 985 1102 990 1103
rect 992 1102 997 1103
rect 473 1003 476 1007
rect 476 1003 477 1007
rect 477 1003 478 1007
rect 480 1003 481 1007
rect 481 1003 482 1007
rect 482 1003 485 1007
rect 473 1002 478 1003
rect 480 1002 485 1003
rect 985 903 988 907
rect 988 903 989 907
rect 989 903 990 907
rect 992 903 993 907
rect 993 903 994 907
rect 994 903 997 907
rect 985 902 990 903
rect 992 902 997 903
rect 473 803 476 807
rect 476 803 477 807
rect 477 803 478 807
rect 480 803 481 807
rect 481 803 482 807
rect 482 803 485 807
rect 473 802 478 803
rect 480 802 485 803
rect 985 703 988 707
rect 988 703 989 707
rect 989 703 990 707
rect 992 703 993 707
rect 993 703 994 707
rect 994 703 997 707
rect 985 702 990 703
rect 992 702 997 703
rect 473 603 476 607
rect 476 603 477 607
rect 477 603 478 607
rect 480 603 481 607
rect 481 603 482 607
rect 482 603 485 607
rect 473 602 478 603
rect 480 602 485 603
rect 985 503 988 507
rect 988 503 989 507
rect 989 503 990 507
rect 992 503 993 507
rect 993 503 994 507
rect 994 503 997 507
rect 985 502 990 503
rect 992 502 997 503
rect 473 403 476 407
rect 476 403 477 407
rect 477 403 478 407
rect 480 403 481 407
rect 481 403 482 407
rect 482 403 485 407
rect 473 402 478 403
rect 480 402 485 403
rect 985 303 988 307
rect 988 303 989 307
rect 989 303 990 307
rect 992 303 993 307
rect 993 303 994 307
rect 994 303 997 307
rect 985 302 990 303
rect 992 302 997 303
rect 473 203 476 207
rect 476 203 477 207
rect 477 203 478 207
rect 480 203 481 207
rect 481 203 482 207
rect 482 203 485 207
rect 473 202 478 203
rect 480 202 485 203
rect 985 103 988 107
rect 988 103 989 107
rect 989 103 990 107
rect 992 103 993 107
rect 993 103 994 107
rect 994 103 997 107
rect 985 102 990 103
rect 992 102 997 103
rect 473 3 476 7
rect 476 3 477 7
rect 477 3 478 7
rect 480 3 481 7
rect 481 3 482 7
rect 482 3 485 7
rect 473 2 478 3
rect 480 2 485 3
<< metal6 >>
rect 472 1207 488 1230
rect 472 1202 473 1207
rect 478 1202 480 1207
rect 485 1202 488 1207
rect 472 1007 488 1202
rect 472 1002 473 1007
rect 478 1002 480 1007
rect 485 1002 488 1007
rect 472 807 488 1002
rect 472 802 473 807
rect 478 802 480 807
rect 485 802 488 807
rect 472 607 488 802
rect 472 602 473 607
rect 478 602 480 607
rect 485 602 488 607
rect 472 407 488 602
rect 472 402 473 407
rect 478 402 480 407
rect 485 402 488 407
rect 472 207 488 402
rect 472 202 473 207
rect 478 202 480 207
rect 485 202 488 207
rect 472 7 488 202
rect 472 2 473 7
rect 478 2 480 7
rect 485 2 488 7
rect 472 -30 488 2
rect 984 1107 1000 1230
rect 984 1102 985 1107
rect 990 1102 992 1107
rect 997 1102 1000 1107
rect 984 907 1000 1102
rect 984 902 985 907
rect 990 902 992 907
rect 997 902 1000 907
rect 984 707 1000 902
rect 984 702 985 707
rect 990 702 992 707
rect 997 702 1000 707
rect 984 507 1000 702
rect 984 502 985 507
rect 990 502 992 507
rect 997 502 1000 507
rect 984 307 1000 502
rect 984 302 985 307
rect 990 302 992 307
rect 997 302 1000 307
rect 984 107 1000 302
rect 984 102 985 107
rect 990 102 992 107
rect 997 102 1000 107
rect 984 -30 1000 102
use DFFPOSX1  DFFPOSX1_10
timestamp 1537539148
transform 1 0 4 0 1 1105
box 0 0 96 100
use INVX1  INVX1_13
timestamp 1537539148
transform 1 0 100 0 1 1105
box 0 0 16 100
use NOR2X1  NOR2X1_25
timestamp 1537539148
transform 1 0 116 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_27
timestamp 1537539148
transform 1 0 140 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_31
timestamp 1537539148
transform 1 0 164 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_25
timestamp 1537539148
transform 1 0 188 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_32
timestamp 1537539148
transform 1 0 212 0 1 1105
box 0 0 24 100
use AOI21X1  AOI21X1_7
timestamp 1537539148
transform 1 0 236 0 1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_17
timestamp 1537539148
transform -1 0 292 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_29
timestamp 1537539148
transform 1 0 292 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_17
timestamp 1537539148
transform 1 0 316 0 1 1105
box 0 0 24 100
use BUFX4  BUFX4_9
timestamp 1537539148
transform -1 0 372 0 1 1105
box 0 0 32 100
use BUFX2  BUFX2_26
timestamp 1537539148
transform 1 0 372 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_30
timestamp 1537539148
transform 1 0 396 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_22
timestamp 1537539148
transform 1 0 420 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_21
timestamp 1537539148
transform 1 0 444 0 1 1105
box 0 0 24 100
use FILL  FILL_11_0_0
timestamp 1537539148
transform 1 0 468 0 1 1105
box 0 0 8 100
use FILL  FILL_11_0_1
timestamp 1537539148
transform 1 0 476 0 1 1105
box 0 0 8 100
use NAND2X1  NAND2X1_6
timestamp 1537539148
transform 1 0 484 0 1 1105
box 0 0 24 100
use INVX2  INVX2_3
timestamp 1537539148
transform -1 0 524 0 1 1105
box 0 0 16 100
use DFFPOSX1  DFFPOSX1_3
timestamp 1537539148
transform 1 0 524 0 1 1105
box 0 0 96 100
use NAND2X1  NAND2X1_7
timestamp 1537539148
transform 1 0 620 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_20
timestamp 1537539148
transform 1 0 644 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_18
timestamp 1537539148
transform 1 0 668 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_19
timestamp 1537539148
transform -1 0 716 0 1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_1
timestamp 1537539148
transform -1 0 748 0 1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_2
timestamp 1537539148
transform 1 0 748 0 1 1105
box 0 0 32 100
use AOI22X1  AOI22X1_1
timestamp 1537539148
transform -1 0 820 0 1 1105
box 0 0 40 100
use INVX2  INVX2_5
timestamp 1537539148
transform -1 0 836 0 1 1105
box 0 0 16 100
use DFFPOSX1  DFFPOSX1_18
timestamp 1537539148
transform 1 0 836 0 1 1105
box 0 0 96 100
use INVX1  INVX1_9
timestamp 1537539148
transform -1 0 948 0 1 1105
box 0 0 16 100
use INVX1  INVX1_12
timestamp 1537539148
transform 1 0 948 0 1 1105
box 0 0 16 100
use AOI21X1  AOI21X1_6
timestamp 1537539148
transform 1 0 964 0 1 1105
box 0 0 32 100
use FILL  FILL_11_1_0
timestamp 1537539148
transform -1 0 1004 0 1 1105
box 0 0 8 100
use FILL  FILL_11_1_1
timestamp 1537539148
transform -1 0 1012 0 1 1105
box 0 0 8 100
use AOI21X1  AOI21X1_1
timestamp 1537539148
transform -1 0 1044 0 1 1105
box 0 0 32 100
use INVX1  INVX1_7
timestamp 1537539148
transform -1 0 1060 0 1 1105
box 0 0 16 100
use NAND2X1  NAND2X1_15
timestamp 1537539148
transform 1 0 1060 0 1 1105
box 0 0 24 100
use NAND2X1  NAND2X1_19
timestamp 1537539148
transform 1 0 1084 0 1 1105
box 0 0 24 100
use NAND2X1  NAND2X1_9
timestamp 1537539148
transform 1 0 1108 0 1 1105
box 0 0 24 100
use NAND2X1  NAND2X1_12
timestamp 1537539148
transform 1 0 1132 0 1 1105
box 0 0 24 100
use INVX1  INVX1_10
timestamp 1537539148
transform 1 0 1156 0 1 1105
box 0 0 16 100
use AOI21X1  AOI21X1_3
timestamp 1537539148
transform 1 0 1172 0 1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_17
timestamp 1537539148
transform -1 0 1228 0 1 1105
box 0 0 24 100
use NAND2X1  NAND2X1_8
timestamp 1537539148
transform -1 0 1252 0 1 1105
box 0 0 24 100
use NAND2X1  NAND2X1_16
timestamp 1537539148
transform 1 0 1252 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_62
timestamp 1537539148
transform -1 0 1300 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_46
timestamp 1537539148
transform 1 0 1300 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_49
timestamp 1537539148
transform 1 0 1324 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_44
timestamp 1537539148
transform 1 0 1348 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_47
timestamp 1537539148
transform 1 0 1372 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_45
timestamp 1537539148
transform 1 0 1396 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_48
timestamp 1537539148
transform 1 0 1420 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_59
timestamp 1537539148
transform 1 0 1444 0 1 1105
box 0 0 24 100
use FILL  FILL_12_1
timestamp 1537539148
transform 1 0 1468 0 1 1105
box 0 0 8 100
use FILL  FILL_12_2
timestamp 1537539148
transform 1 0 1476 0 1 1105
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_16
timestamp 1537539148
transform 1 0 4 0 -1 1105
box 0 0 96 100
use INVX1  INVX1_19
timestamp 1537539148
transform 1 0 100 0 -1 1105
box 0 0 16 100
use NOR2X1  NOR2X1_31
timestamp 1537539148
transform 1 0 116 0 -1 1105
box 0 0 24 100
use BUFX4  BUFX4_13
timestamp 1537539148
transform -1 0 172 0 -1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_29
timestamp 1537539148
transform -1 0 196 0 -1 1105
box 0 0 24 100
use INVX1  INVX1_17
timestamp 1537539148
transform -1 0 212 0 -1 1105
box 0 0 16 100
use DFFPOSX1  DFFPOSX1_2
timestamp 1537539148
transform 1 0 212 0 -1 1105
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_7
timestamp 1537539148
transform 1 0 308 0 -1 1105
box 0 0 96 100
use NOR2X1  NOR2X1_22
timestamp 1537539148
transform -1 0 428 0 -1 1105
box 0 0 24 100
use AOI21X1  AOI21X1_12
timestamp 1537539148
transform -1 0 460 0 -1 1105
box 0 0 32 100
use FILL  FILL_10_0_0
timestamp 1537539148
transform -1 0 468 0 -1 1105
box 0 0 8 100
use FILL  FILL_10_0_1
timestamp 1537539148
transform -1 0 476 0 -1 1105
box 0 0 8 100
use BUFX4  BUFX4_14
timestamp 1537539148
transform -1 0 508 0 -1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_12
timestamp 1537539148
transform 1 0 508 0 -1 1105
box 0 0 24 100
use AOI21X1  AOI21X1_8
timestamp 1537539148
transform 1 0 532 0 -1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_18
timestamp 1537539148
transform -1 0 588 0 -1 1105
box 0 0 24 100
use NOR2X1  NOR2X1_11
timestamp 1537539148
transform -1 0 612 0 -1 1105
box 0 0 24 100
use INVX1  INVX1_4
timestamp 1537539148
transform 1 0 612 0 -1 1105
box 0 0 16 100
use AOI21X1  AOI21X1_9
timestamp 1537539148
transform 1 0 628 0 -1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_19
timestamp 1537539148
transform -1 0 684 0 -1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_4
timestamp 1537539148
transform -1 0 780 0 -1 1105
box 0 0 96 100
use NOR2X1  NOR2X1_13
timestamp 1537539148
transform 1 0 780 0 -1 1105
box 0 0 24 100
use AOI21X1  AOI21X1_2
timestamp 1537539148
transform -1 0 836 0 -1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_29
timestamp 1537539148
transform -1 0 868 0 -1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_28
timestamp 1537539148
transform 1 0 868 0 -1 1105
box 0 0 32 100
use INVX2  INVX2_4
timestamp 1537539148
transform 1 0 900 0 -1 1105
box 0 0 16 100
use OAI21X1  OAI21X1_5
timestamp 1537539148
transform -1 0 948 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_3
timestamp 1537539148
transform 1 0 948 0 -1 1105
box 0 0 32 100
use FILL  FILL_10_1_0
timestamp 1537539148
transform -1 0 988 0 -1 1105
box 0 0 8 100
use FILL  FILL_10_1_1
timestamp 1537539148
transform -1 0 996 0 -1 1105
box 0 0 8 100
use OAI22X1  OAI22X1_1
timestamp 1537539148
transform -1 0 1036 0 -1 1105
box 0 0 40 100
use MUX2X1  MUX2X1_3
timestamp 1537539148
transform 1 0 1036 0 -1 1105
box 0 0 48 100
use OAI21X1  OAI21X1_4
timestamp 1537539148
transform 1 0 1084 0 -1 1105
box 0 0 32 100
use INVX1  INVX1_11
timestamp 1537539148
transform 1 0 1116 0 -1 1105
box 0 0 16 100
use MUX2X1  MUX2X1_1
timestamp 1537539148
transform 1 0 1132 0 -1 1105
box 0 0 48 100
use OAI21X1  OAI21X1_18
timestamp 1537539148
transform -1 0 1212 0 -1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_3
timestamp 1537539148
transform 1 0 1212 0 -1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_17
timestamp 1537539148
transform 1 0 1244 0 -1 1105
box 0 0 32 100
use BUFX4  BUFX4_21
timestamp 1537539148
transform 1 0 1276 0 -1 1105
box 0 0 32 100
use BUFX2  BUFX2_39
timestamp 1537539148
transform -1 0 1332 0 -1 1105
box 0 0 24 100
use BUFX2  BUFX2_67
timestamp 1537539148
transform -1 0 1356 0 -1 1105
box 0 0 24 100
use BUFX2  BUFX2_40
timestamp 1537539148
transform 1 0 1356 0 -1 1105
box 0 0 24 100
use BUFX4  BUFX4_18
timestamp 1537539148
transform 1 0 1380 0 -1 1105
box 0 0 32 100
use BUFX2  BUFX2_42
timestamp 1537539148
transform -1 0 1436 0 -1 1105
box 0 0 24 100
use BUFX2  BUFX2_41
timestamp 1537539148
transform -1 0 1460 0 -1 1105
box 0 0 24 100
use BUFX2  BUFX2_43
timestamp 1537539148
transform 1 0 1460 0 -1 1105
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_17
timestamp 1537539148
transform 1 0 4 0 1 905
box 0 0 96 100
use INVX1  INVX1_20
timestamp 1537539148
transform 1 0 100 0 1 905
box 0 0 16 100
use NOR2X1  NOR2X1_32
timestamp 1537539148
transform 1 0 116 0 1 905
box 0 0 24 100
use BUFX4  BUFX4_16
timestamp 1537539148
transform -1 0 172 0 1 905
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_14
timestamp 1537539148
transform 1 0 172 0 1 905
box 0 0 96 100
use BUFX2  BUFX2_28
timestamp 1537539148
transform 1 0 268 0 1 905
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_15
timestamp 1537539148
transform 1 0 292 0 1 905
box 0 0 96 100
use NOR2X1  NOR2X1_30
timestamp 1537539148
transform -1 0 412 0 1 905
box 0 0 24 100
use INVX1  INVX1_18
timestamp 1537539148
transform -1 0 428 0 1 905
box 0 0 16 100
use NOR2X1  NOR2X1_21
timestamp 1537539148
transform 1 0 428 0 1 905
box 0 0 24 100
use BUFX4  BUFX4_15
timestamp 1537539148
transform -1 0 484 0 1 905
box 0 0 32 100
use FILL  FILL_9_0_0
timestamp 1537539148
transform -1 0 492 0 1 905
box 0 0 8 100
use FILL  FILL_9_0_1
timestamp 1537539148
transform -1 0 500 0 1 905
box 0 0 8 100
use AOI21X1  AOI21X1_11
timestamp 1537539148
transform -1 0 532 0 1 905
box 0 0 32 100
use BUFX4  BUFX4_17
timestamp 1537539148
transform 1 0 532 0 1 905
box 0 0 32 100
use BUFX2  BUFX2_24
timestamp 1537539148
transform 1 0 564 0 1 905
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_9
timestamp 1537539148
transform -1 0 684 0 1 905
box 0 0 96 100
use NOR2X1  NOR2X1_24
timestamp 1537539148
transform 1 0 684 0 1 905
box 0 0 24 100
use AOI21X1  AOI21X1_14
timestamp 1537539148
transform -1 0 740 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_12
timestamp 1537539148
transform 1 0 740 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_13
timestamp 1537539148
transform 1 0 772 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_30
timestamp 1537539148
transform 1 0 804 0 1 905
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_25
timestamp 1537539148
transform 1 0 836 0 1 905
box 0 0 96 100
use OAI21X1  OAI21X1_8
timestamp 1537539148
transform 1 0 932 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_9
timestamp 1537539148
transform 1 0 964 0 1 905
box 0 0 32 100
use FILL  FILL_9_1_0
timestamp 1537539148
transform -1 0 1004 0 1 905
box 0 0 8 100
use FILL  FILL_9_1_1
timestamp 1537539148
transform -1 0 1012 0 1 905
box 0 0 8 100
use MUX2X1  MUX2X1_4
timestamp 1537539148
transform -1 0 1060 0 1 905
box 0 0 48 100
use NOR2X1  NOR2X1_14
timestamp 1537539148
transform -1 0 1084 0 1 905
box 0 0 24 100
use NOR2X1  NOR2X1_9
timestamp 1537539148
transform 1 0 1084 0 1 905
box 0 0 24 100
use XNOR2X1  XNOR2X1_1
timestamp 1537539148
transform -1 0 1164 0 1 905
box 0 0 56 100
use AOI21X1  AOI21X1_4
timestamp 1537539148
transform -1 0 1196 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_22
timestamp 1537539148
transform 1 0 1196 0 1 905
box 0 0 32 100
use INVX1  INVX1_5
timestamp 1537539148
transform -1 0 1244 0 1 905
box 0 0 16 100
use MUX2X1  MUX2X1_2
timestamp 1537539148
transform 1 0 1244 0 1 905
box 0 0 48 100
use BUFX2  BUFX2_36
timestamp 1537539148
transform -1 0 1316 0 1 905
box 0 0 24 100
use BUFX2  BUFX2_37
timestamp 1537539148
transform -1 0 1340 0 1 905
box 0 0 24 100
use BUFX4  BUFX4_22
timestamp 1537539148
transform 1 0 1340 0 1 905
box 0 0 32 100
use BUFX2  BUFX2_35
timestamp 1537539148
transform -1 0 1396 0 1 905
box 0 0 24 100
use BUFX2  BUFX2_38
timestamp 1537539148
transform -1 0 1420 0 1 905
box 0 0 24 100
use BUFX2  BUFX2_68
timestamp 1537539148
transform -1 0 1444 0 1 905
box 0 0 24 100
use BUFX2  BUFX2_63
timestamp 1537539148
transform -1 0 1468 0 1 905
box 0 0 24 100
use FILL  FILL_10_1
timestamp 1537539148
transform 1 0 1468 0 1 905
box 0 0 8 100
use FILL  FILL_10_2
timestamp 1537539148
transform 1 0 1476 0 1 905
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_12
timestamp 1537539148
transform 1 0 4 0 -1 905
box 0 0 96 100
use INVX1  INVX1_15
timestamp 1537539148
transform 1 0 100 0 -1 905
box 0 0 16 100
use NOR2X1  NOR2X1_27
timestamp 1537539148
transform 1 0 116 0 -1 905
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_13
timestamp 1537539148
transform 1 0 140 0 -1 905
box 0 0 96 100
use INVX1  INVX1_16
timestamp 1537539148
transform 1 0 236 0 -1 905
box 0 0 16 100
use NOR2X1  NOR2X1_28
timestamp 1537539148
transform 1 0 252 0 -1 905
box 0 0 24 100
use NOR2X1  NOR2X1_26
timestamp 1537539148
transform -1 0 300 0 -1 905
box 0 0 24 100
use INVX1  INVX1_14
timestamp 1537539148
transform -1 0 316 0 -1 905
box 0 0 16 100
use DFFPOSX1  DFFPOSX1_11
timestamp 1537539148
transform 1 0 316 0 -1 905
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_6
timestamp 1537539148
transform -1 0 508 0 -1 905
box 0 0 96 100
use FILL  FILL_8_0_0
timestamp 1537539148
transform -1 0 516 0 -1 905
box 0 0 8 100
use FILL  FILL_8_0_1
timestamp 1537539148
transform -1 0 524 0 -1 905
box 0 0 8 100
use BUFX4  BUFX4_12
timestamp 1537539148
transform -1 0 556 0 -1 905
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_5
timestamp 1537539148
transform 1 0 556 0 -1 905
box 0 0 96 100
use NOR2X1  NOR2X1_20
timestamp 1537539148
transform 1 0 652 0 -1 905
box 0 0 24 100
use AOI21X1  AOI21X1_10
timestamp 1537539148
transform -1 0 708 0 -1 905
box 0 0 32 100
use INVX1  INVX1_6
timestamp 1537539148
transform 1 0 708 0 -1 905
box 0 0 16 100
use AND2X2  AND2X2_10
timestamp 1537539148
transform 1 0 724 0 -1 905
box 0 0 32 100
use OAI21X1  OAI21X1_27
timestamp 1537539148
transform 1 0 756 0 -1 905
box 0 0 32 100
use INVX2  INVX2_2
timestamp 1537539148
transform -1 0 804 0 -1 905
box 0 0 16 100
use NAND3X1  NAND3X1_2
timestamp 1537539148
transform 1 0 804 0 -1 905
box 0 0 32 100
use AOI21X1  AOI21X1_5
timestamp 1537539148
transform -1 0 868 0 -1 905
box 0 0 32 100
use OAI21X1  OAI21X1_25
timestamp 1537539148
transform -1 0 900 0 -1 905
box 0 0 32 100
use OAI21X1  OAI21X1_20
timestamp 1537539148
transform 1 0 900 0 -1 905
box 0 0 32 100
use NAND3X1  NAND3X1_7
timestamp 1537539148
transform -1 0 964 0 -1 905
box 0 0 32 100
use INVX4  INVX4_2
timestamp 1537539148
transform 1 0 964 0 -1 905
box 0 0 24 100
use FILL  FILL_8_1_0
timestamp 1537539148
transform 1 0 988 0 -1 905
box 0 0 8 100
use FILL  FILL_8_1_1
timestamp 1537539148
transform 1 0 996 0 -1 905
box 0 0 8 100
use BUFX2  BUFX2_55
timestamp 1537539148
transform 1 0 1004 0 -1 905
box 0 0 24 100
use AND2X2  AND2X2_2
timestamp 1537539148
transform -1 0 1060 0 -1 905
box 0 0 32 100
use OAI21X1  OAI21X1_21
timestamp 1537539148
transform 1 0 1060 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_9
timestamp 1537539148
transform 1 0 1092 0 -1 905
box 0 0 32 100
use OAI21X1  OAI21X1_24
timestamp 1537539148
transform 1 0 1124 0 -1 905
box 0 0 32 100
use OAI21X1  OAI21X1_23
timestamp 1537539148
transform -1 0 1188 0 -1 905
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_24
timestamp 1537539148
transform 1 0 1188 0 -1 905
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_19
timestamp 1537539148
transform 1 0 1284 0 -1 905
box 0 0 96 100
use BUFX4  BUFX4_20
timestamp 1537539148
transform -1 0 1412 0 -1 905
box 0 0 32 100
use BUFX2  BUFX2_70
timestamp 1537539148
transform -1 0 1436 0 -1 905
box 0 0 24 100
use BUFX2  BUFX2_75
timestamp 1537539148
transform 1 0 1436 0 -1 905
box 0 0 24 100
use BUFX2  BUFX2_58
timestamp 1537539148
transform -1 0 1484 0 -1 905
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_8
timestamp 1537539148
transform 1 0 4 0 1 705
box 0 0 96 100
use XOR2X1  XOR2X1_1
timestamp 1537539148
transform -1 0 156 0 1 705
box 0 0 56 100
use NOR2X1  NOR2X1_23
timestamp 1537539148
transform -1 0 180 0 1 705
box 0 0 24 100
use AOI21X1  AOI21X1_13
timestamp 1537539148
transform -1 0 212 0 1 705
box 0 0 32 100
use BUFX2  BUFX2_23
timestamp 1537539148
transform 1 0 212 0 1 705
box 0 0 24 100
use BUFX2  BUFX2_69
timestamp 1537539148
transform -1 0 260 0 1 705
box 0 0 24 100
use BUFX2  BUFX2_66
timestamp 1537539148
transform 1 0 260 0 1 705
box 0 0 24 100
use BUFX2  BUFX2_74
timestamp 1537539148
transform 1 0 284 0 1 705
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_22
timestamp 1537539148
transform -1 0 404 0 1 705
box 0 0 96 100
use NOR2X1  NOR2X1_10
timestamp 1537539148
transform 1 0 404 0 1 705
box 0 0 24 100
use NAND3X1  NAND3X1_1
timestamp 1537539148
transform -1 0 460 0 1 705
box 0 0 32 100
use FILL  FILL_7_0_0
timestamp 1537539148
transform 1 0 460 0 1 705
box 0 0 8 100
use FILL  FILL_7_0_1
timestamp 1537539148
transform 1 0 468 0 1 705
box 0 0 8 100
use OAI21X1  OAI21X1_26
timestamp 1537539148
transform 1 0 476 0 1 705
box 0 0 32 100
use NOR2X1  NOR2X1_8
timestamp 1537539148
transform 1 0 508 0 1 705
box 0 0 24 100
use OAI21X1  OAI21X1_14
timestamp 1537539148
transform 1 0 532 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_3
timestamp 1537539148
transform 1 0 564 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_8
timestamp 1537539148
transform -1 0 628 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_5
timestamp 1537539148
transform -1 0 660 0 1 705
box 0 0 32 100
use NOR3X1  NOR3X1_1
timestamp 1537539148
transform -1 0 724 0 1 705
box 0 0 64 100
use NAND2X1  NAND2X1_11
timestamp 1537539148
transform 1 0 724 0 1 705
box 0 0 24 100
use AND2X2  AND2X2_6
timestamp 1537539148
transform 1 0 748 0 1 705
box 0 0 32 100
use NAND2X1  NAND2X1_13
timestamp 1537539148
transform 1 0 780 0 1 705
box 0 0 24 100
use NAND3X1  NAND3X1_4
timestamp 1537539148
transform -1 0 836 0 1 705
box 0 0 32 100
use OAI21X1  OAI21X1_15
timestamp 1537539148
transform 1 0 836 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_6
timestamp 1537539148
transform 1 0 868 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_8
timestamp 1537539148
transform -1 0 932 0 1 705
box 0 0 32 100
use INVX4  INVX4_1
timestamp 1537539148
transform 1 0 932 0 1 705
box 0 0 24 100
use OAI21X1  OAI21X1_16
timestamp 1537539148
transform 1 0 956 0 1 705
box 0 0 32 100
use FILL  FILL_7_1_0
timestamp 1537539148
transform 1 0 988 0 1 705
box 0 0 8 100
use FILL  FILL_7_1_1
timestamp 1537539148
transform 1 0 996 0 1 705
box 0 0 8 100
use AND2X2  AND2X2_7
timestamp 1537539148
transform 1 0 1004 0 1 705
box 0 0 32 100
use OAI21X1  OAI21X1_19
timestamp 1537539148
transform 1 0 1036 0 1 705
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_23
timestamp 1537539148
transform 1 0 1068 0 1 705
box 0 0 96 100
use INVX2  INVX2_1
timestamp 1537539148
transform -1 0 1180 0 1 705
box 0 0 16 100
use BUFX2  BUFX2_56
timestamp 1537539148
transform 1 0 1180 0 1 705
box 0 0 24 100
use BUFX2  BUFX2_52
timestamp 1537539148
transform 1 0 1204 0 1 705
box 0 0 24 100
use XOR2X1  XOR2X1_3
timestamp 1537539148
transform -1 0 1284 0 1 705
box 0 0 56 100
use DFFPOSX1  DFFPOSX1_28
timestamp 1537539148
transform 1 0 1284 0 1 705
box 0 0 96 100
use BUFX2  BUFX2_54
timestamp 1537539148
transform 1 0 1380 0 1 705
box 0 0 24 100
use BUFX2  BUFX2_53
timestamp 1537539148
transform 1 0 1404 0 1 705
box 0 0 24 100
use BUFX2  BUFX2_73
timestamp 1537539148
transform -1 0 1452 0 1 705
box 0 0 24 100
use BUFX2  BUFX2_71
timestamp 1537539148
transform 1 0 1452 0 1 705
box 0 0 24 100
use FILL  FILL_8_1
timestamp 1537539148
transform 1 0 1476 0 1 705
box 0 0 8 100
use BUFX2  BUFX2_16
timestamp 1537539148
transform -1 0 28 0 -1 705
box 0 0 24 100
use BUFX2  BUFX2_33
timestamp 1537539148
transform -1 0 52 0 -1 705
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_27
timestamp 1537539148
transform -1 0 148 0 -1 705
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_26
timestamp 1537539148
transform 1 0 148 0 -1 705
box 0 0 96 100
use XOR2X1  XOR2X1_2
timestamp 1537539148
transform -1 0 300 0 -1 705
box 0 0 56 100
use BUFX2  BUFX2_65
timestamp 1537539148
transform -1 0 324 0 -1 705
box 0 0 24 100
use BUFX2  BUFX2_64
timestamp 1537539148
transform -1 0 348 0 -1 705
box 0 0 24 100
use BUFX2  BUFX2_72
timestamp 1537539148
transform 1 0 348 0 -1 705
box 0 0 24 100
use BUFX4  BUFX4_19
timestamp 1537539148
transform -1 0 404 0 -1 705
box 0 0 32 100
use BUFX2  BUFX2_34
timestamp 1537539148
transform 1 0 404 0 -1 705
box 0 0 24 100
use BUFX4  BUFX4_8
timestamp 1537539148
transform -1 0 460 0 -1 705
box 0 0 32 100
use FILL  FILL_6_0_0
timestamp 1537539148
transform 1 0 460 0 -1 705
box 0 0 8 100
use FILL  FILL_6_0_1
timestamp 1537539148
transform 1 0 468 0 -1 705
box 0 0 8 100
use BUFX4  BUFX4_2
timestamp 1537539148
transform 1 0 476 0 -1 705
box 0 0 32 100
use BUFX2  BUFX2_61
timestamp 1537539148
transform 1 0 508 0 -1 705
box 0 0 24 100
use AND2X2  AND2X2_5
timestamp 1537539148
transform -1 0 564 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_11
timestamp 1537539148
transform -1 0 596 0 -1 705
box 0 0 32 100
use INVX2  INVX2_6
timestamp 1537539148
transform -1 0 612 0 -1 705
box 0 0 16 100
use NOR2X1  NOR2X1_16
timestamp 1537539148
transform 1 0 612 0 -1 705
box 0 0 24 100
use AOI22X1  AOI22X1_2
timestamp 1537539148
transform 1 0 636 0 -1 705
box 0 0 40 100
use INVX1  INVX1_8
timestamp 1537539148
transform -1 0 692 0 -1 705
box 0 0 16 100
use NAND2X1  NAND2X1_10
timestamp 1537539148
transform 1 0 692 0 -1 705
box 0 0 24 100
use OAI21X1  OAI21X1_6
timestamp 1537539148
transform -1 0 748 0 -1 705
box 0 0 32 100
use NOR3X1  NOR3X1_2
timestamp 1537539148
transform 1 0 748 0 -1 705
box 0 0 64 100
use NOR2X1  NOR2X1_15
timestamp 1537539148
transform 1 0 812 0 -1 705
box 0 0 24 100
use NAND2X1  NAND2X1_14
timestamp 1537539148
transform 1 0 836 0 -1 705
box 0 0 24 100
use NOR3X1  NOR3X1_3
timestamp 1537539148
transform 1 0 860 0 -1 705
box 0 0 64 100
use NAND2X1  NAND2X1_18
timestamp 1537539148
transform -1 0 948 0 -1 705
box 0 0 24 100
use BUFX4  BUFX4_5
timestamp 1537539148
transform 1 0 948 0 -1 705
box 0 0 32 100
use FILL  FILL_6_1_0
timestamp 1537539148
transform 1 0 980 0 -1 705
box 0 0 8 100
use FILL  FILL_6_1_1
timestamp 1537539148
transform 1 0 988 0 -1 705
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_20
timestamp 1537539148
transform 1 0 996 0 -1 705
box 0 0 96 100
use NOR2X1  NOR2X1_33
timestamp 1537539148
transform 1 0 1092 0 -1 705
box 0 0 24 100
use INVX1  INVX1_21
timestamp 1537539148
transform -1 0 1132 0 -1 705
box 0 0 16 100
use NOR2X1  NOR2X1_34
timestamp 1537539148
transform 1 0 1132 0 -1 705
box 0 0 24 100
use OAI21X1  OAI21X1_31
timestamp 1537539148
transform 1 0 1156 0 -1 705
box 0 0 32 100
use XNOR2X1  XNOR2X1_2
timestamp 1537539148
transform 1 0 1188 0 -1 705
box 0 0 56 100
use DFFPOSX1  DFFPOSX1_29
timestamp 1537539148
transform 1 0 1244 0 -1 705
box 0 0 96 100
use BUFX2  BUFX2_2
timestamp 1537539148
transform 1 0 1340 0 -1 705
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_1
timestamp 1537539148
transform 1 0 1364 0 -1 705
box 0 0 96 100
use FILL  FILL_7_1
timestamp 1537539148
transform -1 0 1468 0 -1 705
box 0 0 8 100
use FILL  FILL_7_2
timestamp 1537539148
transform -1 0 1476 0 -1 705
box 0 0 8 100
use FILL  FILL_7_3
timestamp 1537539148
transform -1 0 1484 0 -1 705
box 0 0 8 100
use BUFX2  BUFX2_50
timestamp 1537539148
transform -1 0 28 0 1 505
box 0 0 24 100
use BUFX2  BUFX2_51
timestamp 1537539148
transform -1 0 52 0 1 505
box 0 0 24 100
use NOR2X1  NOR2X1_5
timestamp 1537539148
transform 1 0 52 0 1 505
box 0 0 24 100
use NOR2X1  NOR2X1_6
timestamp 1537539148
transform 1 0 76 0 1 505
box 0 0 24 100
use NAND2X1  NAND2X1_4
timestamp 1537539148
transform -1 0 124 0 1 505
box 0 0 24 100
use OR2X2  OR2X2_1
timestamp 1537539148
transform -1 0 156 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_16
timestamp 1537539148
transform 1 0 156 0 1 505
box 0 0 32 100
use INVX1  INVX1_36
timestamp 1537539148
transform 1 0 188 0 1 505
box 0 0 16 100
use AOI21X1  AOI21X1_26
timestamp 1537539148
transform 1 0 204 0 1 505
box 0 0 32 100
use NOR2X1  NOR2X1_59
timestamp 1537539148
transform -1 0 260 0 1 505
box 0 0 24 100
use NAND3X1  NAND3X1_25
timestamp 1537539148
transform -1 0 292 0 1 505
box 0 0 32 100
use INVX1  INVX1_3
timestamp 1537539148
transform 1 0 292 0 1 505
box 0 0 16 100
use NAND2X1  NAND2X1_5
timestamp 1537539148
transform -1 0 332 0 1 505
box 0 0 24 100
use NOR2X1  NOR2X1_7
timestamp 1537539148
transform -1 0 356 0 1 505
box 0 0 24 100
use NOR2X1  NOR2X1_1
timestamp 1537539148
transform 1 0 356 0 1 505
box 0 0 24 100
use NAND2X1  NAND2X1_1
timestamp 1537539148
transform 1 0 380 0 1 505
box 0 0 24 100
use INVX1  INVX1_1
timestamp 1537539148
transform -1 0 420 0 1 505
box 0 0 16 100
use BUFX4  BUFX4_4
timestamp 1537539148
transform -1 0 452 0 1 505
box 0 0 32 100
use NOR2X1  NOR2X1_2
timestamp 1537539148
transform 1 0 452 0 1 505
box 0 0 24 100
use FILL  FILL_5_0_0
timestamp 1537539148
transform -1 0 484 0 1 505
box 0 0 8 100
use FILL  FILL_5_0_1
timestamp 1537539148
transform -1 0 492 0 1 505
box 0 0 8 100
use NOR2X1  NOR2X1_4
timestamp 1537539148
transform -1 0 516 0 1 505
box 0 0 24 100
use DFFPOSX1  DFFPOSX1_21
timestamp 1537539148
transform -1 0 612 0 1 505
box 0 0 96 100
use OAI21X1  OAI21X1_7
timestamp 1537539148
transform -1 0 644 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_4
timestamp 1537539148
transform 1 0 644 0 1 505
box 0 0 32 100
use OAI21X1  OAI21X1_10
timestamp 1537539148
transform 1 0 676 0 1 505
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_35
timestamp 1537539148
transform 1 0 708 0 1 505
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_31
timestamp 1537539148
transform 1 0 804 0 1 505
box 0 0 96 100
use NOR3X1  NOR3X1_4
timestamp 1537539148
transform -1 0 964 0 1 505
box 0 0 64 100
use AND2X2  AND2X2_11
timestamp 1537539148
transform 1 0 964 0 1 505
box 0 0 32 100
use FILL  FILL_5_1_0
timestamp 1537539148
transform 1 0 996 0 1 505
box 0 0 8 100
use FILL  FILL_5_1_1
timestamp 1537539148
transform 1 0 1004 0 1 505
box 0 0 8 100
use NAND2X1  NAND2X1_20
timestamp 1537539148
transform 1 0 1012 0 1 505
box 0 0 24 100
use INVX2  INVX2_7
timestamp 1537539148
transform 1 0 1036 0 1 505
box 0 0 16 100
use OR2X2  OR2X2_2
timestamp 1537539148
transform 1 0 1052 0 1 505
box 0 0 32 100
use NAND2X1  NAND2X1_21
timestamp 1537539148
transform -1 0 1108 0 1 505
box 0 0 24 100
use AND2X2  AND2X2_12
timestamp 1537539148
transform -1 0 1140 0 1 505
box 0 0 32 100
use NAND3X1  NAND3X1_9
timestamp 1537539148
transform -1 0 1172 0 1 505
box 0 0 32 100
use OAI21X1  OAI21X1_32
timestamp 1537539148
transform -1 0 1204 0 1 505
box 0 0 32 100
use XNOR2X1  XNOR2X1_3
timestamp 1537539148
transform 1 0 1204 0 1 505
box 0 0 56 100
use DFFPOSX1  DFFPOSX1_30
timestamp 1537539148
transform 1 0 1260 0 1 505
box 0 0 96 100
use BUFX2  BUFX2_3
timestamp 1537539148
transform 1 0 1356 0 1 505
box 0 0 24 100
use BUFX2  BUFX2_1
timestamp 1537539148
transform 1 0 1380 0 1 505
box 0 0 24 100
use BUFX2  BUFX2_4
timestamp 1537539148
transform 1 0 1404 0 1 505
box 0 0 24 100
use BUFX2  BUFX2_5
timestamp 1537539148
transform 1 0 1428 0 1 505
box 0 0 24 100
use BUFX2  BUFX2_57
timestamp 1537539148
transform -1 0 1476 0 1 505
box 0 0 24 100
use FILL  FILL_6_1
timestamp 1537539148
transform 1 0 1476 0 1 505
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_44
timestamp 1537539148
transform 1 0 4 0 -1 505
box 0 0 96 100
use NAND2X1  NAND2X1_36
timestamp 1537539148
transform -1 0 124 0 -1 505
box 0 0 24 100
use NOR2X1  NOR2X1_45
timestamp 1537539148
transform 1 0 124 0 -1 505
box 0 0 24 100
use NAND2X1  NAND2X1_33
timestamp 1537539148
transform 1 0 148 0 -1 505
box 0 0 24 100
use NAND3X1  NAND3X1_18
timestamp 1537539148
transform -1 0 204 0 -1 505
box 0 0 32 100
use NAND3X1  NAND3X1_17
timestamp 1537539148
transform -1 0 236 0 -1 505
box 0 0 32 100
use OAI21X1  OAI21X1_49
timestamp 1537539148
transform -1 0 268 0 -1 505
box 0 0 32 100
use INVX2  INVX2_10
timestamp 1537539148
transform -1 0 284 0 -1 505
box 0 0 16 100
use NOR3X1  NOR3X1_12
timestamp 1537539148
transform -1 0 348 0 -1 505
box 0 0 64 100
use OR2X2  OR2X2_4
timestamp 1537539148
transform 1 0 348 0 -1 505
box 0 0 32 100
use NOR2X1  NOR2X1_49
timestamp 1537539148
transform -1 0 404 0 -1 505
box 0 0 24 100
use OAI21X1  OAI21X1_58
timestamp 1537539148
transform 1 0 404 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_37
timestamp 1537539148
transform -1 0 460 0 -1 505
box 0 0 24 100
use NAND2X1  NAND2X1_2
timestamp 1537539148
transform 1 0 460 0 -1 505
box 0 0 24 100
use FILL  FILL_4_0_0
timestamp 1537539148
transform -1 0 492 0 -1 505
box 0 0 8 100
use FILL  FILL_4_0_1
timestamp 1537539148
transform -1 0 500 0 -1 505
box 0 0 8 100
use INVX1  INVX1_2
timestamp 1537539148
transform -1 0 516 0 -1 505
box 0 0 16 100
use NAND2X1  NAND2X1_3
timestamp 1537539148
transform -1 0 540 0 -1 505
box 0 0 24 100
use NOR2X1  NOR2X1_3
timestamp 1537539148
transform 1 0 540 0 -1 505
box 0 0 24 100
use AND2X2  AND2X2_1
timestamp 1537539148
transform 1 0 564 0 -1 505
box 0 0 32 100
use BUFX4  BUFX4_7
timestamp 1537539148
transform 1 0 596 0 -1 505
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_36
timestamp 1537539148
transform 1 0 628 0 -1 505
box 0 0 96 100
use BUFX4  BUFX4_11
timestamp 1537539148
transform 1 0 724 0 -1 505
box 0 0 32 100
use BUFX4  BUFX4_1
timestamp 1537539148
transform 1 0 756 0 -1 505
box 0 0 32 100
use INVX8  INVX8_1
timestamp 1537539148
transform -1 0 828 0 -1 505
box 0 0 40 100
use DFFPOSX1  DFFPOSX1_33
timestamp 1537539148
transform 1 0 828 0 -1 505
box 0 0 96 100
use XNOR2X1  XNOR2X1_6
timestamp 1537539148
transform -1 0 980 0 -1 505
box 0 0 56 100
use FILL  FILL_4_1_0
timestamp 1537539148
transform 1 0 980 0 -1 505
box 0 0 8 100
use FILL  FILL_4_1_1
timestamp 1537539148
transform 1 0 988 0 -1 505
box 0 0 8 100
use XNOR2X1  XNOR2X1_4
timestamp 1537539148
transform 1 0 996 0 -1 505
box 0 0 56 100
use AOI21X1  AOI21X1_15
timestamp 1537539148
transform 1 0 1052 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_23
timestamp 1537539148
transform -1 0 1108 0 -1 505
box 0 0 24 100
use OAI21X1  OAI21X1_33
timestamp 1537539148
transform -1 0 1140 0 -1 505
box 0 0 32 100
use OAI21X1  OAI21X1_35
timestamp 1537539148
transform -1 0 1172 0 -1 505
box 0 0 32 100
use NAND3X1  NAND3X1_11
timestamp 1537539148
transform 1 0 1172 0 -1 505
box 0 0 32 100
use NAND3X1  NAND3X1_10
timestamp 1537539148
transform -1 0 1236 0 -1 505
box 0 0 32 100
use OAI21X1  OAI21X1_34
timestamp 1537539148
transform -1 0 1268 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_22
timestamp 1537539148
transform 1 0 1268 0 -1 505
box 0 0 24 100
use INVX1  INVX1_22
timestamp 1537539148
transform -1 0 1308 0 -1 505
box 0 0 16 100
use XNOR2X1  XNOR2X1_5
timestamp 1537539148
transform 1 0 1308 0 -1 505
box 0 0 56 100
use DFFPOSX1  DFFPOSX1_32
timestamp 1537539148
transform 1 0 1364 0 -1 505
box 0 0 96 100
use FILL  FILL_5_1
timestamp 1537539148
transform -1 0 1468 0 -1 505
box 0 0 8 100
use FILL  FILL_5_2
timestamp 1537539148
transform -1 0 1476 0 -1 505
box 0 0 8 100
use FILL  FILL_5_3
timestamp 1537539148
transform -1 0 1484 0 -1 505
box 0 0 8 100
use NOR3X1  NOR3X1_18
timestamp 1537539148
transform -1 0 68 0 1 305
box 0 0 64 100
use NOR2X1  NOR2X1_55
timestamp 1537539148
transform 1 0 68 0 1 305
box 0 0 24 100
use INVX1  INVX1_32
timestamp 1537539148
transform 1 0 92 0 1 305
box 0 0 16 100
use NAND3X1  NAND3X1_19
timestamp 1537539148
transform -1 0 140 0 1 305
box 0 0 32 100
use NAND2X1  NAND2X1_32
timestamp 1537539148
transform -1 0 164 0 1 305
box 0 0 24 100
use NAND2X1  NAND2X1_38
timestamp 1537539148
transform 1 0 164 0 1 305
box 0 0 24 100
use OAI21X1  OAI21X1_50
timestamp 1537539148
transform 1 0 188 0 1 305
box 0 0 32 100
use NOR2X1  NOR2X1_51
timestamp 1537539148
transform -1 0 244 0 1 305
box 0 0 24 100
use NOR2X1  NOR2X1_50
timestamp 1537539148
transform -1 0 268 0 1 305
box 0 0 24 100
use NOR2X1  NOR2X1_60
timestamp 1537539148
transform -1 0 292 0 1 305
box 0 0 24 100
use NOR3X1  NOR3X1_14
timestamp 1537539148
transform 1 0 292 0 1 305
box 0 0 64 100
use INVX4  INVX4_4
timestamp 1537539148
transform 1 0 356 0 1 305
box 0 0 24 100
use NAND3X1  NAND3X1_20
timestamp 1537539148
transform -1 0 412 0 1 305
box 0 0 32 100
use INVX1  INVX1_37
timestamp 1537539148
transform 1 0 412 0 1 305
box 0 0 16 100
use OAI21X1  OAI21X1_59
timestamp 1537539148
transform -1 0 460 0 1 305
box 0 0 32 100
use FILL  FILL_3_0_0
timestamp 1537539148
transform 1 0 460 0 1 305
box 0 0 8 100
use FILL  FILL_3_0_1
timestamp 1537539148
transform 1 0 468 0 1 305
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_43
timestamp 1537539148
transform 1 0 476 0 1 305
box 0 0 96 100
use NAND2X1  NAND2X1_42
timestamp 1537539148
transform 1 0 572 0 1 305
box 0 0 24 100
use NOR2X1  NOR2X1_48
timestamp 1537539148
transform 1 0 596 0 1 305
box 0 0 24 100
use NAND3X1  NAND3X1_16
timestamp 1537539148
transform 1 0 620 0 1 305
box 0 0 32 100
use NOR2X1  NOR2X1_47
timestamp 1537539148
transform -1 0 676 0 1 305
box 0 0 24 100
use OAI21X1  OAI21X1_57
timestamp 1537539148
transform -1 0 708 0 1 305
box 0 0 32 100
use NAND2X1  NAND2X1_43
timestamp 1537539148
transform -1 0 732 0 1 305
box 0 0 24 100
use BUFX4  BUFX4_10
timestamp 1537539148
transform 1 0 732 0 1 305
box 0 0 32 100
use BUFX4  BUFX4_3
timestamp 1537539148
transform 1 0 764 0 1 305
box 0 0 32 100
use XNOR2X1  XNOR2X1_8
timestamp 1537539148
transform -1 0 852 0 1 305
box 0 0 56 100
use XNOR2X1  XNOR2X1_9
timestamp 1537539148
transform -1 0 908 0 1 305
box 0 0 56 100
use BUFX4  BUFX4_6
timestamp 1537539148
transform 1 0 908 0 1 305
box 0 0 32 100
use INVX1  INVX1_24
timestamp 1537539148
transform 1 0 940 0 1 305
box 0 0 16 100
use AND2X2  AND2X2_13
timestamp 1537539148
transform -1 0 988 0 1 305
box 0 0 32 100
use FILL  FILL_3_1_0
timestamp 1537539148
transform 1 0 988 0 1 305
box 0 0 8 100
use FILL  FILL_3_1_1
timestamp 1537539148
transform 1 0 996 0 1 305
box 0 0 8 100
use OAI21X1  OAI21X1_37
timestamp 1537539148
transform 1 0 1004 0 1 305
box 0 0 32 100
use AOI21X1  AOI21X1_18
timestamp 1537539148
transform 1 0 1036 0 1 305
box 0 0 32 100
use AOI21X1  AOI21X1_16
timestamp 1537539148
transform 1 0 1068 0 1 305
box 0 0 32 100
use OAI21X1  OAI21X1_36
timestamp 1537539148
transform 1 0 1100 0 1 305
box 0 0 32 100
use NAND2X1  NAND2X1_25
timestamp 1537539148
transform 1 0 1132 0 1 305
box 0 0 24 100
use AOI21X1  AOI21X1_17
timestamp 1537539148
transform -1 0 1188 0 1 305
box 0 0 32 100
use INVX1  INVX1_23
timestamp 1537539148
transform -1 0 1204 0 1 305
box 0 0 16 100
use NAND2X1  NAND2X1_26
timestamp 1537539148
transform -1 0 1228 0 1 305
box 0 0 24 100
use NOR2X1  NOR2X1_35
timestamp 1537539148
transform -1 0 1252 0 1 305
box 0 0 24 100
use XNOR2X1  XNOR2X1_7
timestamp 1537539148
transform 1 0 1252 0 1 305
box 0 0 56 100
use NAND2X1  NAND2X1_27
timestamp 1537539148
transform -1 0 1332 0 1 305
box 0 0 24 100
use NAND2X1  NAND2X1_24
timestamp 1537539148
transform -1 0 1356 0 1 305
box 0 0 24 100
use BUFX2  BUFX2_11
timestamp 1537539148
transform 1 0 1356 0 1 305
box 0 0 24 100
use BUFX2  BUFX2_9
timestamp 1537539148
transform 1 0 1380 0 1 305
box 0 0 24 100
use BUFX2  BUFX2_7
timestamp 1537539148
transform 1 0 1404 0 1 305
box 0 0 24 100
use BUFX2  BUFX2_6
timestamp 1537539148
transform 1 0 1428 0 1 305
box 0 0 24 100
use BUFX2  BUFX2_60
timestamp 1537539148
transform -1 0 1476 0 1 305
box 0 0 24 100
use FILL  FILL_4_1
timestamp 1537539148
transform 1 0 1476 0 1 305
box 0 0 8 100
use DFFPOSX1  DFFPOSX1_45
timestamp 1537539148
transform 1 0 4 0 -1 305
box 0 0 96 100
use AND2X2  AND2X2_15
timestamp 1537539148
transform 1 0 100 0 -1 305
box 0 0 32 100
use NAND2X1  NAND2X1_41
timestamp 1537539148
transform -1 0 156 0 -1 305
box 0 0 24 100
use INVX1  INVX1_35
timestamp 1537539148
transform -1 0 172 0 -1 305
box 0 0 16 100
use NAND2X1  NAND2X1_39
timestamp 1537539148
transform -1 0 196 0 -1 305
box 0 0 24 100
use NOR2X1  NOR2X1_42
timestamp 1537539148
transform 1 0 196 0 -1 305
box 0 0 24 100
use OAI21X1  OAI21X1_46
timestamp 1537539148
transform -1 0 252 0 -1 305
box 0 0 32 100
use OAI22X1  OAI22X1_4
timestamp 1537539148
transform 1 0 252 0 -1 305
box 0 0 40 100
use INVX1  INVX1_34
timestamp 1537539148
transform 1 0 292 0 -1 305
box 0 0 16 100
use INVX4  INVX4_3
timestamp 1537539148
transform -1 0 332 0 -1 305
box 0 0 24 100
use NAND2X1  NAND2X1_44
timestamp 1537539148
transform -1 0 356 0 -1 305
box 0 0 24 100
use INVX1  INVX1_31
timestamp 1537539148
transform 1 0 356 0 -1 305
box 0 0 16 100
use OAI21X1  OAI21X1_47
timestamp 1537539148
transform 1 0 372 0 -1 305
box 0 0 32 100
use NOR3X1  NOR3X1_11
timestamp 1537539148
transform -1 0 468 0 -1 305
box 0 0 64 100
use FILL  FILL_2_0_0
timestamp 1537539148
transform 1 0 468 0 -1 305
box 0 0 8 100
use FILL  FILL_2_0_1
timestamp 1537539148
transform 1 0 476 0 -1 305
box 0 0 8 100
use OAI21X1  OAI21X1_52
timestamp 1537539148
transform 1 0 484 0 -1 305
box 0 0 32 100
use OAI21X1  OAI21X1_53
timestamp 1537539148
transform -1 0 548 0 -1 305
box 0 0 32 100
use INVX2  INVX2_11
timestamp 1537539148
transform -1 0 564 0 -1 305
box 0 0 16 100
use NOR3X1  NOR3X1_10
timestamp 1537539148
transform -1 0 628 0 -1 305
box 0 0 64 100
use DFFPOSX1  DFFPOSX1_46
timestamp 1537539148
transform 1 0 628 0 -1 305
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_41
timestamp 1537539148
transform 1 0 724 0 -1 305
box 0 0 96 100
use INVX1  INVX1_28
timestamp 1537539148
transform 1 0 820 0 -1 305
box 0 0 16 100
use XNOR2X1  XNOR2X1_13
timestamp 1537539148
transform -1 0 892 0 -1 305
box 0 0 56 100
use OAI21X1  OAI21X1_44
timestamp 1537539148
transform 1 0 892 0 -1 305
box 0 0 32 100
use AOI21X1  AOI21X1_22
timestamp 1537539148
transform -1 0 956 0 -1 305
box 0 0 32 100
use OAI21X1  OAI21X1_38
timestamp 1537539148
transform 1 0 956 0 -1 305
box 0 0 32 100
use FILL  FILL_2_1_0
timestamp 1537539148
transform 1 0 988 0 -1 305
box 0 0 8 100
use FILL  FILL_2_1_1
timestamp 1537539148
transform 1 0 996 0 -1 305
box 0 0 8 100
use BUFX2  BUFX2_14
timestamp 1537539148
transform 1 0 1004 0 -1 305
box 0 0 24 100
use BUFX2  BUFX2_12
timestamp 1537539148
transform 1 0 1028 0 -1 305
box 0 0 24 100
use NAND3X1  NAND3X1_12
timestamp 1537539148
transform 1 0 1052 0 -1 305
box 0 0 32 100
use INVX1  INVX1_25
timestamp 1537539148
transform -1 0 1100 0 -1 305
box 0 0 16 100
use OAI21X1  OAI21X1_39
timestamp 1537539148
transform 1 0 1100 0 -1 305
box 0 0 32 100
use NOR2X1  NOR2X1_38
timestamp 1537539148
transform 1 0 1132 0 -1 305
box 0 0 24 100
use NOR2X1  NOR2X1_37
timestamp 1537539148
transform 1 0 1156 0 -1 305
box 0 0 24 100
use NAND3X1  NAND3X1_13
timestamp 1537539148
transform 1 0 1180 0 -1 305
box 0 0 32 100
use NOR3X1  NOR3X1_5
timestamp 1537539148
transform 1 0 1212 0 -1 305
box 0 0 64 100
use NOR2X1  NOR2X1_36
timestamp 1537539148
transform 1 0 1276 0 -1 305
box 0 0 24 100
use OR2X2  OR2X2_3
timestamp 1537539148
transform -1 0 1332 0 -1 305
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_34
timestamp 1537539148
transform 1 0 1332 0 -1 305
box 0 0 96 100
use BUFX2  BUFX2_10
timestamp 1537539148
transform 1 0 1428 0 -1 305
box 0 0 24 100
use BUFX2  BUFX2_8
timestamp 1537539148
transform -1 0 1476 0 -1 305
box 0 0 24 100
use FILL  FILL_3_1
timestamp 1537539148
transform -1 0 1484 0 -1 305
box 0 0 8 100
use NAND3X1  NAND3X1_23
timestamp 1537539148
transform -1 0 36 0 1 105
box 0 0 32 100
use NOR3X1  NOR3X1_19
timestamp 1537539148
transform 1 0 36 0 1 105
box 0 0 64 100
use OAI21X1  OAI21X1_55
timestamp 1537539148
transform -1 0 132 0 1 105
box 0 0 32 100
use OAI21X1  OAI21X1_54
timestamp 1537539148
transform -1 0 164 0 1 105
box 0 0 32 100
use NAND3X1  NAND3X1_21
timestamp 1537539148
transform 1 0 164 0 1 105
box 0 0 32 100
use OAI21X1  OAI21X1_51
timestamp 1537539148
transform 1 0 196 0 1 105
box 0 0 32 100
use OAI22X1  OAI22X1_3
timestamp 1537539148
transform -1 0 268 0 1 105
box 0 0 40 100
use NOR2X1  NOR2X1_43
timestamp 1537539148
transform -1 0 292 0 1 105
box 0 0 24 100
use AOI21X1  AOI21X1_25
timestamp 1537539148
transform 1 0 292 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_58
timestamp 1537539148
transform 1 0 324 0 1 105
box 0 0 24 100
use NOR2X1  NOR2X1_44
timestamp 1537539148
transform 1 0 348 0 1 105
box 0 0 24 100
use OAI21X1  OAI21X1_56
timestamp 1537539148
transform 1 0 372 0 1 105
box 0 0 32 100
use INVX1  INVX1_30
timestamp 1537539148
transform -1 0 420 0 1 105
box 0 0 16 100
use NAND2X1  NAND2X1_31
timestamp 1537539148
transform 1 0 420 0 1 105
box 0 0 24 100
use NAND3X1  NAND3X1_22
timestamp 1537539148
transform 1 0 444 0 1 105
box 0 0 32 100
use FILL  FILL_1_0_0
timestamp 1537539148
transform -1 0 484 0 1 105
box 0 0 8 100
use FILL  FILL_1_0_1
timestamp 1537539148
transform -1 0 492 0 1 105
box 0 0 8 100
use NAND2X1  NAND2X1_34
timestamp 1537539148
transform -1 0 516 0 1 105
box 0 0 24 100
use OAI22X1  OAI22X1_2
timestamp 1537539148
transform -1 0 556 0 1 105
box 0 0 40 100
use NAND3X1  NAND3X1_15
timestamp 1537539148
transform 1 0 556 0 1 105
box 0 0 32 100
use NAND3X1  NAND3X1_24
timestamp 1537539148
transform 1 0 588 0 1 105
box 0 0 32 100
use NOR3X1  NOR3X1_9
timestamp 1537539148
transform 1 0 620 0 1 105
box 0 0 64 100
use NAND2X1  NAND2X1_35
timestamp 1537539148
transform -1 0 708 0 1 105
box 0 0 24 100
use NOR3X1  NOR3X1_13
timestamp 1537539148
transform 1 0 708 0 1 105
box 0 0 64 100
use DFFPOSX1  DFFPOSX1_39
timestamp 1537539148
transform 1 0 772 0 1 105
box 0 0 96 100
use NAND2X1  NAND2X1_29
timestamp 1537539148
transform 1 0 868 0 1 105
box 0 0 24 100
use NOR3X1  NOR3X1_8
timestamp 1537539148
transform 1 0 892 0 1 105
box 0 0 64 100
use NAND3X1  NAND3X1_14
timestamp 1537539148
transform -1 0 988 0 1 105
box 0 0 32 100
use FILL  FILL_1_1_0
timestamp 1537539148
transform -1 0 996 0 1 105
box 0 0 8 100
use FILL  FILL_1_1_1
timestamp 1537539148
transform -1 0 1004 0 1 105
box 0 0 8 100
use OAI21X1  OAI21X1_43
timestamp 1537539148
transform -1 0 1036 0 1 105
box 0 0 32 100
use INVX1  INVX1_29
timestamp 1537539148
transform 1 0 1036 0 1 105
box 0 0 16 100
use OAI21X1  OAI21X1_45
timestamp 1537539148
transform -1 0 1084 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_41
timestamp 1537539148
transform -1 0 1108 0 1 105
box 0 0 24 100
use NOR3X1  NOR3X1_7
timestamp 1537539148
transform 1 0 1108 0 1 105
box 0 0 64 100
use AOI21X1  AOI21X1_20
timestamp 1537539148
transform 1 0 1172 0 1 105
box 0 0 32 100
use AOI21X1  AOI21X1_19
timestamp 1537539148
transform 1 0 1204 0 1 105
box 0 0 32 100
use INVX2  INVX2_8
timestamp 1537539148
transform -1 0 1252 0 1 105
box 0 0 16 100
use XOR2X1  XOR2X1_4
timestamp 1537539148
transform 1 0 1252 0 1 105
box 0 0 56 100
use XOR2X1  XOR2X1_5
timestamp 1537539148
transform 1 0 1308 0 1 105
box 0 0 56 100
use DFFPOSX1  DFFPOSX1_42
timestamp 1537539148
transform 1 0 1364 0 1 105
box 0 0 96 100
use FILL  FILL_2_1
timestamp 1537539148
transform 1 0 1460 0 1 105
box 0 0 8 100
use FILL  FILL_2_2
timestamp 1537539148
transform 1 0 1468 0 1 105
box 0 0 8 100
use FILL  FILL_2_3
timestamp 1537539148
transform 1 0 1476 0 1 105
box 0 0 8 100
use NOR3X1  NOR3X1_17
timestamp 1537539148
transform -1 0 68 0 -1 105
box 0 0 64 100
use NOR2X1  NOR2X1_54
timestamp 1537539148
transform 1 0 68 0 -1 105
box 0 0 24 100
use AOI21X1  AOI21X1_23
timestamp 1537539148
transform 1 0 92 0 -1 105
box 0 0 32 100
use NOR2X1  NOR2X1_52
timestamp 1537539148
transform -1 0 148 0 -1 105
box 0 0 24 100
use NOR3X1  NOR3X1_15
timestamp 1537539148
transform -1 0 212 0 -1 105
box 0 0 64 100
use INVX2  INVX2_13
timestamp 1537539148
transform -1 0 228 0 -1 105
box 0 0 16 100
use NAND2X1  NAND2X1_40
timestamp 1537539148
transform 1 0 228 0 -1 105
box 0 0 24 100
use OAI21X1  OAI21X1_48
timestamp 1537539148
transform -1 0 284 0 -1 105
box 0 0 32 100
use INVX1  INVX1_33
timestamp 1537539148
transform -1 0 300 0 -1 105
box 0 0 16 100
use NOR3X1  NOR3X1_16
timestamp 1537539148
transform 1 0 300 0 -1 105
box 0 0 64 100
use NOR2X1  NOR2X1_53
timestamp 1537539148
transform -1 0 388 0 -1 105
box 0 0 24 100
use NOR3X1  NOR3X1_20
timestamp 1537539148
transform 1 0 388 0 -1 105
box 0 0 64 100
use NOR2X1  NOR2X1_57
timestamp 1537539148
transform -1 0 476 0 -1 105
box 0 0 24 100
use FILL  FILL_0_0_0
timestamp 1537539148
transform 1 0 476 0 -1 105
box 0 0 8 100
use FILL  FILL_0_0_1
timestamp 1537539148
transform 1 0 484 0 -1 105
box 0 0 8 100
use NOR2X1  NOR2X1_46
timestamp 1537539148
transform 1 0 492 0 -1 105
box 0 0 24 100
use INVX2  INVX2_12
timestamp 1537539148
transform 1 0 516 0 -1 105
box 0 0 16 100
use NOR2X1  NOR2X1_56
timestamp 1537539148
transform -1 0 556 0 -1 105
box 0 0 24 100
use AOI21X1  AOI21X1_24
timestamp 1537539148
transform 1 0 556 0 -1 105
box 0 0 32 100
use DFFPOSX1  DFFPOSX1_40
timestamp 1537539148
transform -1 0 684 0 -1 105
box 0 0 96 100
use XNOR2X1  XNOR2X1_11
timestamp 1537539148
transform 1 0 684 0 -1 105
box 0 0 56 100
use INVX2  INVX2_9
timestamp 1537539148
transform 1 0 740 0 -1 105
box 0 0 16 100
use XNOR2X1  XNOR2X1_12
timestamp 1537539148
transform -1 0 812 0 -1 105
box 0 0 56 100
use NAND2X1  NAND2X1_28
timestamp 1537539148
transform -1 0 836 0 -1 105
box 0 0 24 100
use NOR2X1  NOR2X1_40
timestamp 1537539148
transform 1 0 836 0 -1 105
box 0 0 24 100
use NAND2X1  NAND2X1_30
timestamp 1537539148
transform -1 0 884 0 -1 105
box 0 0 24 100
use INVX1  INVX1_27
timestamp 1537539148
transform 1 0 884 0 -1 105
box 0 0 16 100
use AOI21X1  AOI21X1_21
timestamp 1537539148
transform 1 0 900 0 -1 105
box 0 0 32 100
use OAI21X1  OAI21X1_42
timestamp 1537539148
transform 1 0 932 0 -1 105
box 0 0 32 100
use AND2X2  AND2X2_14
timestamp 1537539148
transform -1 0 996 0 -1 105
box 0 0 32 100
use FILL  FILL_0_1_0
timestamp 1537539148
transform -1 0 1004 0 -1 105
box 0 0 8 100
use FILL  FILL_0_1_1
timestamp 1537539148
transform -1 0 1012 0 -1 105
box 0 0 8 100
use NOR3X1  NOR3X1_6
timestamp 1537539148
transform -1 0 1076 0 -1 105
box 0 0 64 100
use OAI21X1  OAI21X1_41
timestamp 1537539148
transform -1 0 1108 0 -1 105
box 0 0 32 100
use INVX1  INVX1_26
timestamp 1537539148
transform -1 0 1124 0 -1 105
box 0 0 16 100
use NOR2X1  NOR2X1_39
timestamp 1537539148
transform -1 0 1148 0 -1 105
box 0 0 24 100
use OAI21X1  OAI21X1_40
timestamp 1537539148
transform 1 0 1148 0 -1 105
box 0 0 32 100
use XNOR2X1  XNOR2X1_10
timestamp 1537539148
transform 1 0 1180 0 -1 105
box 0 0 56 100
use DFFPOSX1  DFFPOSX1_38
timestamp 1537539148
transform 1 0 1236 0 -1 105
box 0 0 96 100
use DFFPOSX1  DFFPOSX1_37
timestamp 1537539148
transform 1 0 1332 0 -1 105
box 0 0 96 100
use BUFX2  BUFX2_13
timestamp 1537539148
transform 1 0 1428 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_15
timestamp 1537539148
transform -1 0 1476 0 -1 105
box 0 0 24 100
use FILL  FILL_1_1
timestamp 1537539148
transform -1 0 1484 0 -1 105
box 0 0 8 100
<< labels >>
rlabel metal6 s 472 -30 488 -22 8 vdd
port 0 nsew
rlabel metal6 s 984 -30 1000 -22 8 gnd
port 1 nsew
rlabel metal2 s 352 1230 352 1230 6 clk
port 2 nsew
rlabel metal2 s 1024 1230 1024 1230 6 INPD<0>
port 3 nsew
rlabel metal2 s 984 1230 984 1230 6 INPD<1>
port 4 nsew
rlabel metal2 s 968 1230 968 1230 6 INPD<2>
port 5 nsew
rlabel metal2 s 944 1230 944 1230 6 INPD<3>
port 6 nsew
rlabel metal2 s 928 1230 928 1230 6 INPD<4>
port 7 nsew
rlabel metal2 s 904 1230 904 1230 6 INPD<5>
port 8 nsew
rlabel metal2 s 888 1230 888 1230 6 INPD<6>
port 9 nsew
rlabel metal2 s 864 1230 864 1230 6 INPD<7>
port 10 nsew
rlabel metal2 s 848 1230 848 1230 6 INPD<8>
port 11 nsew
rlabel metal2 s 824 1230 824 1230 6 INPD<9>
port 12 nsew
rlabel metal2 s 808 1230 808 1230 6 INPD<10>
port 13 nsew
rlabel metal2 s 784 1230 784 1230 6 INPD<11>
port 14 nsew
rlabel metal2 s 768 1230 768 1230 6 INPD<12>
port 15 nsew
rlabel metal2 s 744 1230 744 1230 6 INPD<13>
port 16 nsew
rlabel metal2 s 728 1230 728 1230 6 INPD<14>
port 17 nsew
rlabel metal2 s 704 1230 704 1230 6 INPD<15>
port 18 nsew
rlabel metal2 s 1040 1230 1040 1230 6 RDATA<0>
port 19 nsew
rlabel metal2 s 1064 1230 1064 1230 6 RDATA<1>
port 20 nsew
rlabel metal2 s 1080 1230 1080 1230 6 RDATA<2>
port 21 nsew
rlabel metal2 s 1104 1230 1104 1230 6 RDATA<3>
port 22 nsew
rlabel metal2 s 1120 1230 1120 1230 6 RDATA<4>
port 23 nsew
rlabel metal2 s 1144 1230 1144 1230 6 RDATA<5>
port 24 nsew
rlabel metal2 s 1160 1230 1160 1230 6 RDATA<6>
port 25 nsew
rlabel metal2 s 1184 1230 1184 1230 6 RDATA<7>
port 26 nsew
rlabel metal2 s 560 -20 560 -20 8 RF
port 27 nsew
rlabel metal2 s 520 -20 520 -20 8 WF
port 28 nsew
rlabel metal2 s 272 -20 272 -20 8 NEXTOP<0>
port 29 nsew
rlabel metal2 s 232 -20 232 -20 8 NEXTOP<1>
port 30 nsew
rlabel metal2 s 72 -20 72 -20 8 NEXTOP<2>
port 31 nsew
rlabel metal3 s -24 680 -24 680 4 IR
port 32 nsew
rlabel metal3 s -24 660 -24 660 4 OW
port 33 nsew
rlabel metal2 s 688 1230 688 1230 6 OUTPD<0>
port 34 nsew
rlabel metal2 s 664 1230 664 1230 6 OUTPD<1>
port 35 nsew
rlabel metal2 s 648 1230 648 1230 6 OUTPD<2>
port 36 nsew
rlabel metal2 s 624 1230 624 1230 6 OUTPD<3>
port 37 nsew
rlabel metal2 s 608 1230 608 1230 6 OUTPD<4>
port 38 nsew
rlabel metal2 s 584 1230 584 1230 6 OUTPD<5>
port 39 nsew
rlabel metal2 s 568 1230 568 1230 6 OUTPD<6>
port 40 nsew
rlabel metal2 s 544 1230 544 1230 6 OUTPD<7>
port 41 nsew
rlabel metal2 s 528 1230 528 1230 6 OUTPD<8>
port 42 nsew
rlabel metal2 s 488 1230 488 1230 6 OUTPD<9>
port 43 nsew
rlabel metal2 s 472 1230 472 1230 6 OUTPD<10>
port 44 nsew
rlabel metal2 s 448 1230 448 1230 6 OUTPD<11>
port 45 nsew
rlabel metal2 s 432 1230 432 1230 6 OUTPD<12>
port 46 nsew
rlabel metal2 s 408 1230 408 1230 6 OUTPD<13>
port 47 nsew
rlabel metal2 s 392 1230 392 1230 6 OUTPD<14>
port 48 nsew
rlabel metal2 s 368 1230 368 1230 6 OUTPD<15>
port 49 nsew
rlabel metal3 s 1512 360 1512 360 6 reset
port 50 nsew
rlabel metal3 s -24 580 -24 580 4 RD
port 51 nsew
rlabel metal3 s -24 560 -24 560 4 WD
port 52 nsew
rlabel metal3 s 1512 760 1512 760 6 WDATA<0>
port 53 nsew
rlabel metal3 s 1512 780 1512 780 6 WDATA<1>
port 54 nsew
rlabel metal3 s 1512 800 1512 800 6 WDATA<2>
port 55 nsew
rlabel metal3 s 1512 860 1512 860 6 WDATA<3>
port 56 nsew
rlabel metal3 s 1512 880 1512 880 6 WDATA<4>
port 57 nsew
rlabel metal3 s 1512 900 1512 900 6 WDATA<5>
port 58 nsew
rlabel metal3 s 1512 920 1512 920 6 WDATA<6>
port 59 nsew
rlabel metal3 s 1512 1060 1512 1060 6 WDATA<7>
port 60 nsew
rlabel metal3 s 1512 680 1512 680 6 DP<0>
port 61 nsew
rlabel metal3 s 1512 660 1512 660 6 DP<1>
port 62 nsew
rlabel metal3 s 1512 620 1512 620 6 DP<2>
port 63 nsew
rlabel metal3 s 1512 600 1512 600 6 DP<3>
port 64 nsew
rlabel metal3 s 1512 580 1512 580 6 DP<4>
port 65 nsew
rlabel metal3 s 1512 560 1512 560 6 DP<5>
port 66 nsew
rlabel metal3 s 1512 540 1512 540 6 DP<6>
port 67 nsew
rlabel metal3 s 1512 520 1512 520 6 DP<7>
port 68 nsew
rlabel metal3 s 1512 500 1512 500 6 DP<8>
port 69 nsew
rlabel metal3 s 1512 480 1512 480 6 DP<9>
port 70 nsew
rlabel metal3 s 1512 460 1512 460 6 DP<10>
port 71 nsew
rlabel metal3 s 1512 440 1512 440 6 DP<11>
port 72 nsew
rlabel metal3 s 1512 420 1512 420 6 DP<12>
port 73 nsew
rlabel metal3 s 1512 400 1512 400 6 DP<13>
port 74 nsew
rlabel metal3 s 1512 380 1512 380 6 DP<14>
port 75 nsew
rlabel metal2 s 1200 1230 1200 1230 6 PCDELTA<0>
port 76 nsew
rlabel metal2 s 1224 1230 1224 1230 6 PCDELTA<1>
port 77 nsew
rlabel metal2 s 1240 1230 1240 1230 6 PCDELTA<2>
port 78 nsew
rlabel metal2 s 1264 1230 1264 1230 6 PCDELTA<3>
port 79 nsew
rlabel metal2 s 1280 1230 1280 1230 6 PCDELTA<4>
port 80 nsew
rlabel metal2 s 1304 1230 1304 1230 6 PCDELTA<5>
port 81 nsew
rlabel metal2 s 1320 1230 1320 1230 6 PCDELTA<6>
port 82 nsew
rlabel metal2 s 1344 1230 1344 1230 6 PCDELTA<7>
port 83 nsew
rlabel metal2 s 1360 1230 1360 1230 6 PCDELTA<8>
port 84 nsew
rlabel metal2 s 1384 1230 1384 1230 6 PCDELTA<9>
port 85 nsew
rlabel metal2 s 1400 1230 1400 1230 6 PCDELTA<10>
port 86 nsew
rlabel metal2 s 1424 1230 1424 1230 6 PCDELTA<11>
port 87 nsew
rlabel metal2 s 1440 1230 1440 1230 6 PCDELTA<12>
port 88 nsew
rlabel metal2 s 1464 1230 1464 1230 6 PCDELTA<13>
port 89 nsew
rlabel metal2 s 1480 1230 1480 1230 6 PCDELTA<14>
port 90 nsew
rlabel metal2 s 1504 1230 1504 1230 6 PCDELTA<15>
port 91 nsew
<< end >>
